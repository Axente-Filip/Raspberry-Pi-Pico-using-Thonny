PK   �M�Z�
Bv;	  �I     cirkitFile.json͛mo�8ǿ��{sXY>�R�]��� �m�z/� D��U����6[���Pv����f^\P!��!E�����ר��|�*�ί>�nS�Mt��2����lǥl��fշ��]�G�_�s�?�}\���M��S$��q��.V&1����J	f��4lŢ�w������'�8���5N���'Oq��;$w	G�Ǒ�q${	G�Ǒ�q$ɟ��{H��?��O �H��?��O ��H�$�?��x��I$ɟD�'��I$ɟB�����al��"v�e�g&Ne)��W2�	��gN���{?K����ؙ%?:��#g��t�̒���Y��a3K~:j�a3`��|m�v��+�~"TF�E�x�$^�M�%!�bH��$^2�ॡ����i��4 s�9�aN1��X�P,��`�ł�bAC���X�P,h(4K�%Œ�(AC���X�P,i(�4K�%Ŋ�bEC��H��L����W���x��s�X/�rnNK��bH��p	�\������sڻ�m�io�}gkdڋ�"H�H/�ċ&�x1$^R/uD����i��4�r�9��aN�0����P,h(Dk0ł�bAC���X�P,h(4�%Œ�bIt���X�P,i(�4K�%Œ�bEC���X]�xvڋ�r�f��x/�rvڋ�r1(g��x/Crvڋ�r1 秽On �m��~�Y�r_�o�~�:�Y�k[x������v.�L�h?��6�x5۹m����s[��!��V�g��6F/�z��+�^#�	Ro���ϰ���ȱr,�!�Rȱr,�"ǒ(�$
�Z�%Q`IX�D�%Q`IX�D�%QbI��mK�Ē(�$J,�K�Ē(�$*,�
K�:C��,�?��3K��L ��&1�3a4;�������?B�3�U�����x܄�mN@B��i9\.	��KÕ�e�J��B��b��CU��P���<T�>"(��;(DP��A!�B�
2(dPȡ;A!�B�
2(dP��PA!����/�:|�z����ahW�/c�K����6�5����*�uy�5d�e���M�K�O[3����ʾE��v��ô>���+0l��j>@?���u}��6<��a�0;ۦ�6"��ܷ�_57�6�.m��`���m�����:�Ƕ꼋��n��l�-m�o;ߝk\�#���:�]��x]t'|!��T����VWY&2�L�J�Мg����[FeR���<.�4�3fҸ�B�%��wZK3�v����?�^FR�m���Y���ڮ/v��h������~r�I&��R���r��b,�fT���(}.��Z�zz�'��Wf?X��&��b��\��i�J*_���;�N��,r'���&5���$U��}+:������j��}[�:�4�D�F�o��}����ذbf������H�&��MGFdl����rd&��D��	��ɶ&\M,cǆ	����HlL�G�jb?��8�'�q���&��LfW�\���=��c�a�qa��Z-˶v�[~�����.�|�}q-��%�(
�	X�J�sE��,��<U6+X����u��F������iYb�,6���Y'>�i��B2ŬWYY�A�頿��Vkm|��Hc�����J�(����f��Gb#�+sh���L�=,�Eac�9�0'�vf�����w\��1�{�~���澪��s��&EK�X���2&N�byɘ`i6��um�j훑%l��<���z�gq愌��e)t^*=��n7~ܛF�;��F$��8eY�L���%l���|Y����;*��?x&���7��}��C����*�A>���'c�����\�7���ے/��˲����@4FL{����F��y�:�cmR��,���b�e"0��10��X���/�!����38��!F�k89��&:p��̌�{�$� H�)L!�H�g��yĊ��]����b�����[|��k��~Z@s��v��,�P{q�;�\���6��'�P�}���m{�σ��#n:�����~;�����}�����d�h�~�3�~_;�)�8�	,��?��>V��~��p̊����@
����o1��N�|߬m���mC~�հgaOq���*I
X���y��X��H]����YG�YYԌ#�V�+�CZ��{3*O�����~����P>�������ތ�ӧ�K�����6n��oaF"�wĆ���e�4���,UC���r�=�I�^�D�����}�(%T7~�N�8�2w[�{����|�?�����Or��bUׯʗ�]\�X>7�C��w/�;[�hn{�V[HL�+t�!V������	���PK   �M�Z��'S4  N4  /   images/90a7334e-e219-40c9-b800-02625da96495.pngN4�ˉPNG

   IHDR   d   h    U/   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  3�IDATx�՝`TU��ϴL	%	B�RBQDD@PAAt��]W�ow-k��������.������ ,�(�HCK }f��w^f2̤�=�̔w߼w�=�ν��y}�e!y�y����Ȏ�"n�T��r��IO���پ�U���Ex�+��ꒂ�~ԯ8�ׁ���'�g�24(`�q����M7%��/����~�j���7"۶�С�RV��^pɹ�64���U�u���>�<�%K
䤓h�r��}=K_������C�����P���1��#��>[��~�U��}�z����*��S_l%����)�����r�2.O��Ehs�U"��f���K$��< )�{�G�:�'�|ⓑ#E
E��'�[n�T��>�m]����\�˂��ϊL��"~(r�i�^`����w�RC�)I�+)y����/�H�7u�]tQ����_�Zz����x��1�)Y�� �{.�O�0O\!�QHGap�2�ԫ�ݧ��|0A����rs��MS%wđ��{;)i�,neH���3}��_�Zd�J�7�E�"2]��~��g�L�${�5���ɦ�m�S���r�ؘ'��ʕ�K׊J�Ȍb��r���׋�%��ײ3;S��l�m��l��6���i�d���0��_���B��C�B�r�"���*�f)/^%e��I�<|��y��$}����AM�|�m��ms�r�h���F2\a���I;�ح����r�$U�kG�]w��=y�l��Z�^>J�5I�j뗟z���<K�N�'2d�a�a�����od]����'JQjJE��d��Y��l/�&|#=f,�mg���^;rUfH�֪vv��q]q�U۪w9��f�\���uf��:?��d���#���j�X��E��U�//)��$��T<e����4m���	��z�u�4ٶK��Y*��EZ�����C�8m?�]�h�v�x��|��9cI��;U����ޤ���Ų�yS���F���J���v������.�y}3�<ִ�^�Ld�Jt�����B�kSC]����V$���/\|�K�}���DJZ���\^��)�$oks�/Ido�a�b@wّ�!��2I�[�������'�HMBu��;+�S��'!��϶mi����9����0#%��������WJqj�4[��mUe�ʒ=�'���ڰ�JK����F3��{�O�;>�|�V٧����-�3��*���f��h����[����5޾���H<ʰ�u���̿�z��>�3�Zm:��Q�v�v�]�����֠���������F�	O x��Mdw����)����.���+̽��W�M��Lc�z}�@U�)_�K^���S^��&i;�M;e�l�������>��ʧ�%�~��G���]��\���H~Jp3^G)aD��c��ztУs�SC�>�kӔ+G�8�Ù2��O��ڭ����xХg�x�%���S5�v��>EM��S�/_^r�� uܮ%���Ǩ��T��Vܮ�/>qC;p�-���W�6RC[�W�g$�!$�,�g\[US˻�\"�j�ν�M�|���p�>�ܽ�/O�s�^I9p�
WP]>��GA���z���J=.�#IjF�K�>a�^��F��_ =� �@:R���Y�ʭT��:������v�9�J�<o�aV�ޢA|�Uu�*����{�P:��Q�g%��׵���~+�+6HA�4i�#P�~�+Ru������T][}�j���w�M��G<G޼�rq����>K��l>���)c�E�1�|�H���'#�$���>��ǋz���uݕ��A�]tT5Q���v����y���Mõ��iW��mX+��ue�g���t��s��~���9cI��U��u�W�@��+�d���m\'z�SI�t]|�Ꮮ��7����f�w������#���[P��f�z�֡%���Ϳ]1NU�mH٤s����|�}�S�Ҷ����|˵������J]��Z�����#��v����U�t���U#���su��� ]]��(_E�b�ۈ�w�x�2w�,;&G�A+�=�I��{��g5_�-[�{B��u#G|6׺�x:]��L�(ݿ]"����3�HR���/������j��i�0l�n�!\���E>�Lr��5�t�:�&y�kOR�����U��AHtʾ"9��y������d��d�"��|�:;S�����,_��N�Ih�t	�{���Q�^����BP�N������v����qr«���+O��[bo�h�w�V^�zA%ṙߪ$�9�0"g��l�%i>���hۓ%�u3u�<=U�Dzz/��d�{_I��r��϶���(��;��pm���08��õ��)�S���d��S%'�%&�F��A��ɹ�B7%������G��89�T���G�h&�gN�[��e���8����9U��կ��N��x%����������M�Vظ����������l���s�nӱ��j����O�X��~��s�$H�����E�Tm�y��W_�6Kտx�-Ӷ��=����v�����3�r�&ӶQ��~��,�S3��^ޭ)3�ϋb
b���':}����'�������*�ʡ�����+]ճ�2U<���YZj1�I��=�i�[�U�}w�0ԣ��K��/��~P�Q>��I�Z8��=��N8�(�&p�Oi۔7ސ#�3���=�3�#n�UjA/W��Ԏb��uj���o�X���"C��w�k�ӻ�ȬY"�9C*PW)�����k�z�Caڢn�f@�!�%\^�P�[/�R[��!/�l�+��{�~���]Wq?^�5��m~��p��2#!�A�bmP�8�U����֎�SN���  ���T��!��O���E´}�]�6����c���� �����w�?�Q�&k���qHaU�e�~5���J���ܟ����ϷG]H��u��S�Q�<��K%b��EE	>�b���F��
ud���99��L��$���)�s�鑢Gi=�L�D?_��Pr���C�f�I֎�z�	��I�L�X�j讦M�F��ok����#���.���{PZ�pÆ6��li�)�vY���E:����w"���wb2�\;F2k�B�)K��ɭ+*�3���Cکc�<S7k&֬Q�����-UQH�s��T9�s�ۨ��"7�j�u+;u����[�~�=�XÀ-�E�{��\T�e\`��1�[�Z#c�Ҭ��2Eǫ�^�l���i��D��p�az4K�]��h��#.���e�ʕ2WGd����*�25�}�3/�Ni�7k��b�ug���L��) ���m ��z��VZ�p�۷i����"���߽[�c��.���JDÑ�����o��'�.����tr�O�_[)���U�Zن�����+�b}]���3�����=�O���6P�ɱ�+:�Ѽv�uIQ[�Ԓ�8{���,�ϛgU��W��,��G�������[����ز���q����ë)Sb�A�1���+{Y!UؒB�}ڹ�ʌ*%D�ߞ�/e:BC����k�F�������ٳ�]p��;����E�`'�tQ)5m�
��kF}-Zd����1U��0������N��)y�7��x�����~��!ne���� ɪ���_W5�4��X;���'���Ƌ:A}�mkG9L@
���	`�3��Ad�+=��I�E�Er0�0
&a����^ƍo��cGP"�H)�*(�_�4j}Hy�� �1qԟz2A��VEB6��m��תD;kL�y}�"����6P�>`��QiT�`G ��/������u���5v���m�
;�"ˆq��ʜ�����%+IH6Y�(��$0Bq�.���ܥ�_��(�����������TC��!lO�J����c�u���Eb���L�]���Pm��|�B��mڈ4h`;�N ģ�;CR ?Q_��g�`�O?��������:��m���_z�h���ۋ�}\(�]�xaHP��zU����Xv�z0�jT��v�T�j+���N'�qHuPxG�����8�(�}��ѣ#��r�Ɉ�p���@0,ր;9���erc� [F�5�����y�tIʔ�ډw�q�	����vh{eƸq�L����V�3JQS{�X�[�H�O%�*E:� ������&(������y �xg��
T��U�z��;w�w�쀽�(J���^ԔG;+SUL��:2�2��*�ڵ����h;��.+��C��c)�$� VQw�R����
��f� o����F�ac8o�bk�p�(�s�xªĸ���Х�7|�C��U�-sn�0]N�Bl0o^�hO��\����UM0"���0<�RS-�LPZvB�ۀ��C�*3ĥ���/�9�#	�^�����j����:���"lN �G���8�K(hZ 	��"i�E�U}�Qo֭j�����1�Օ�Pf��M�o~#5�ATƯA0��AAG�4!ym2L%c��ظ]RH��~c�ȌrnXR��w(�l�B��]@':��%5�����wRO��d���#�`u���T�d42�#�u���?�J��a
�B��ӯ\��eigޡ�/�{R2����<1��=r3.���n��2ȯ2c�cd����έR�.�^�����ǽ1�N����K/�C���wu�7v�zMk�-S��uq��*Z�4�z�F�I�.:��=���󛪦����#M����l{RIٽ�>�}߽<�wW�?�i�����۬,�,��`<��0⎷H:�[���g0���A�9�{�f��F�`�:+�)ʨk����i���Z��X=Ēj����9q�)WW�{��a����yꯒJK��l�5vwV�wHJ�뙗�f�[:���x��ʑÔ!.�7�#�L0�lr7����s:�x
��7�!i �Hy{�U�|l�(����i*�!�0��!H@u�;1�ɝ�Z3��ð�̜2��Ч[���n��ʹ&��}k=e����[�l,LrK�(fTbA'� %��N��2��5�r>$Ź�0LЋt8S<jH�� t��
�"�zC��UJ�~�Qo�T�_T�ڕe��k��n��:�9"�\7V�|��2w��MoD��s�2sn��<-�@�t<���H����ib?#0F����b]s�D��؃�ū"���؅��\�M���m��b�W���x%��lmfڮ�oޔ��;.X���CV޴KG�	�����Շ�Ke}JA���?L`�"p�((4%3�H�����7�(���g�1��������B���1��U�$�];���O�׀�j�!���$S�oG:�����6��������.�z=�o���A5���Q���!�� �y�> ���܇�� NM���#6�#�FB�����|������AOsP��_�`H�`�۷Kd]�Φ�X�Ӱ2���2�r�P�H�������wJ8�[P���.� O�~ء�^�6*X���Y�+���k03��>�tC�HtC�b'3W�r�C��!�OA}_xA������2����.L�����N��~�[Sů�E��Wk+��*1ք%�G�4I;R���QO �H��n-s�IPC�1���2$���5�#��ƨ�q�I��K�$PU�JG�{��qaHc���v�߾{�*Y���"t ���l��إ��A�PjB����6#Y��ʫ���=;/2ꋀ0y_�d��(m�!�jܩ̸3<��X��� �0��%��·HE�R3��D�S�gr���P� 9�l��.��OQ�D_���xT�\	�8С���<С܄��g�-e��E�mS�V�܊����I�֭r���!tFM��ո����^g�?���At�m��'1d���j�*^�q1P�k����">r�HRAΟ|���&�O��!�H�� S�!zQ�zA���C�H��uŸkA��6Ht':��;ࡩ��B��z�z^ \�ZSڨ7]���O��P�HP��CZ�}w��H����C0�R,N�0�OPHu��"�ﶌ�am�. ��b05���abx�ð���$�3��mn�ru��!O��"G��I��5:�߾����+O�R�[p"9��6�TJOY�:�] ��-�fʶ�d= R��$�\L�+3�`17N!"F��a�������36��3�C�4'�C���ڃ�!5�� jp�YDgϞ�_��e���OwC��xA���n�_�7wn]ȥن;�8���.V��o��k&'�DN���ڱɨ+�����Hk��߬�l6$����Z�Y�7� �%ވ�6�B�:�S�>��m�sË���Y!�n)"�]�j�h�@H !���3�]Ed��;��?xV-`�Xb��c�	��%�$�x����H Q1./*
=}�)f���cɏCz��l��T�.����_IՐH��@����tFz�&@:bk���7��E{RHu�.�\�ũ}�9��?C<:��̞-)F��%~����7��a�'�m�,/>�$���]�v����������ˤ���#�Q�0���tp/�^3/Q��4@���-{����g?ϕWZ��@uL�~�|'�L}��\9k�?C�:BW���L�����KU6�Cd���[�����/�d��[��b����O+�g�96G���#�𺯤�uV�&�ܬ��B_iy'���>à�r����Iߩ�z��=X��P��T#��Q�1�������!!{U�e3��v˫���#)�_Q�d2��6Έu ����u�vfn�y�Ζ�칮-]�,����s^O����Ioe��v��{4@�*r��/�����F=�[a>�9mQ��[$4�"Z߀�]�fC�N8$)������M][����'d�19��i�H�����s�w�T��#�����kO��";���-���=Q��g1��{$Z]��f`蝲W
	"��p��ϯ�qXcu���xT s�{E�9�ɬ�R����  ���0�%�c6�@��Bq.5�M�t09�?�}&j%�,�j����QY� ]'�J��j��w�A���x�5�����fU�#�Wl���W��{�1f���s�5Y6��9vE��Ҡ$P� B�K�?�Z*-)�C�3Ɉ8W��Q�Ǆ�Py	>�-bb���i�\�)s�)�;/�f\�gG1���K�6P�+�z
4Ps�C�˓_��J�v`�ݏ�SNuL<�ym�M��ܢ�<�uZqT�>o�Z,��	r"�����0/�ы� 9��b@@qE��yQ)C ���N|EpJ\BD4�(�"e@����p��j�3���h��yq�z,��^�ٸ����\��?�7��� 𑂲�4�_��'���^��S���� �! u�-A� �8� �*AJ�!�C)EZ��M8S��	48������Q�@+�bT#�A{щ���?0����B�� I�ޭ����g�B�&���/����j4��9U�F�f��!k��Ԇ�t战��6�n��:�i��A�]��9 �0x��'O��_�Cᥥŝ��8G����S��n��H
�A�8:�������T�7Rwq�g� $Iv˖Ҡa�T�h���a���l�˨U��V��8S��Z"�;������t�j3.t�`t�E����?�f�Ċ��Y$�Ij���q�$�}�(��Ƕ�s�v)r �WH���D9�ed��s�7�L�F�S$|I���[�!���^�w�OQw���{�Q�T<�f3j4�&��� ��]@I;�,��A˱SHTT�Te����va�W��)�w|�XRC�����L�:
�=�µ�Y��W	+ѣ:��$a�xvw�e K�^�vK�h`���� �ߏ��h2�;�*J�)�J:ϙ�m�-������ŻC�QW�`����a3�K�'������ ���dˈ.QSNnQ���2=Z��q:�<�9�ո�iG�j�*W�j����	�Cg��D�?����uw5	��3��?�q/c	�M���4'ʉ�h�=$ˈ��y%xJ��S1���w�'Յ��L��`�^�*�8ho��	�$z*s"	ё���w�y\9��2�%�ؚH	�xYY�c� T
�Yߩ�X��h��K��M���($)A��t.�!�M�$���GE�C��0�JҶ���Lh�L�Tu¨!��r��b=x)u��pG�l��������ȁ�-@���������ȁ����t��:���M��r�h'��Kҋx�$Yu�ř����ˀiH#5�vڕ�M������e@,��5c���'��`/��X� u0OXBr�6qqQ���1�=T7v��u_C� `a��!X��V'p��Ã�����n��Y׫��9�_7(�w��,�*��d��<������eI���kl*��s+&�c��3H�SQB<Ј���Au�3��H� H�i�=RK����V�}�C�!�
�@8�!F!�_T�1�g��&�Y+�4lP�t��%)~JI�]|�K���5��^w��}:I?e�7���>�6/���=e�TE����瞱���xO�ɴ�h\:��ˉ��/�ޞ����.)2�c�.m��׮@��>m�������|{�q��#ז�]�P?V9-J�HZ<Ƀ��
l$3�q���A{���7�3����x��s�ZPe��Vׯ+a��+F�B(�ح��J��s��%���Fl�ꅱ��Q�������M2K�.�]#�-l}a $ʛ̹�I�R�Li��M7ف��@+KPʽ��Z%��C�u ��n�@6�r�\��T�͆G��G�3��ɱ�_F'���
��@|�r��x�(���e�����y��e:����+7=��̄��K׳�Fu�/ �m��G�k�*`��[^x�B��<+*	I�m�l�SG�0�N����6G��i�.աp�V� ���@o�).TN�G/:v�l~�aq9��6ۧ�X�G�k���?*�QF''P���_ړŋ!*�"F �f	��.��};S����EӉj��0��<�ck��;��bn;'V"�W�Ԓ!< +Q6�(T)�������RM���ԃ +Z�#�0��@5�Q�Au�r� �� 瞩���z8+;v4#h�����JF#��d�>���i��`@B{vK��Ȗ��R2�Ƣ��!�|͒M�*������>O�<�I9͕O��T�#d<��B�6�.K2 8�\�W��T��
w����e+�~�B;�E^�|�:so8�Nӑ�P;b�l}б�g�ĺ�k�/���O%�(�P��UAA����~���w�O��Сr��Y���@؁'?�N�f-�QӢM'�3p(��+�n�y��������fD� 7sŮ�WP@�ix�2�Н á�gْ�zM��ٳw�2�D��تD�G,13�N~���Uu-��zD(��?K
��G3 �8T�Nn�;��ϡ�)�񆥋�Lu�7�\G|w�o���3�)P}��C8�[�ԘgG/��/ji\R�?���8���A	�����L��K�0��L��'_p�K@����S��3�BAf@�C ��d�]Jl������tF<�|?��3���6����DM9�@����:�!�Px
@(� &��}T���[%#�7�xQ�'����	1�`L ���v����D��ɬ�Sjn�5E�u�p�#��{Y}T��@����JW�ty�N�.W��䨕]���Q�*��G���������+
*K��3����/K���ب��0����U��<��lf�Ue\��K�OG�G�E-T��sȉ����Er��E���D,��>��΢wP�D����H�E�ɒ�%P��_6�6zLF���z�9Jm��b�5�Y~���tR� �]��(��%~��VY~��~<+mGI3�ȡ�]ӑ(�|C4�d$�Y.���|F4C�@�#�{�~���#��b2`c�G�����8��K���Cb�$ة�2�QQ���8!�`Y����I���,^3��v��|��m���7�Q271ٳk��߰^�EŒ6���Ę���AB0�n�b�&�7������D\cg��*�F�R��Q���Q�ݫ7!��b@��.a���X��T񐠟�l $��ߠ��8Um��ْ3X�*����]�U�)�W()O=��!0���q}ԍ3�:Xb�h"�J�l�E���F���y���&앪(b��1L�'�KiJ��[����x����=�a�	��$�-��%��{Tz"�D��T�e��'!�V�Fڈ3�
f�B�V�<� G*���x_N*��IE:�)fyvnf۽��
�C(�����l:}��n ��_�RZ����E]�Y9������1��.xV@���T�g�׉U?�j��0���ؒnh��k�g>�EHp46����܃E�`�S��%qpqQ��G%:�Wʁ��'�?bdCT��1�)����F#��	�N�����(�ː���Ee1�)�c^wx��
8��PPP�C%�l"���~�k=(����`�T�=�"���r��`��êb	"p(Z�دHI���pV]8��m]��()�z�<w=2�`�:��CH�\P�v���A}l�n��a����(a)J��}�jcIꢘ�Q�^��jcI"r�����xK�.��@uI�w��2w��ՆSAB��%)¨�d#�:
2�kۼ�D_$fȠ�v�՟�W��*�TD�� B��|xx��J���֫0-z�U����Ԫ����>����@PP@�n0��M(ls�'�֫,S��W	�X%mM-kU*(J%�$m���ю
�9�[o�ls�?��͉���pA9psb[g%�҄�!
�M�91��.>t>6�6D��&ܜ��1�W��T�m�9pbn\�D_��"n��3&Ȧ-��s��R����> C/�EZ�����ۡL���>)�yo�M��d��@g�n�_�~ZJR�oߍ��ˍ{3�"���~�-=?�l�M�{I�dSZ��Y9l�#Qux�H�[U���3ej+%1�U�[�!M��=����.{�vO��
v�òkk7��ۺ�6��IAzZ��f2�0m{����af��3Y����u�4��J���>���m�d�Q�d�{_I���E-op�`��Q��U'h���r@w��Ti#a
�BD�h�H���Űjʔ����$���ڹ�q]:\ܬZf��<𓪬����ܮA���:��s�� m�ݨ+�q˴�Ff0��-��,��l��uB��u�8{��i�d���)~�8QJ��d�'ˎV��WB�����!i�񸇕���/.i;$[�
1�OA�ږ�����]��^[�m���AE�)��%'ɘ�&HL!va@�|����nR���쪘�r$j�"�5�g�)k)5�Ŭ�o/�/*��}�ꋖ�c��&��f������'�;��(}�z/�m��ʣ��	30#y_�;��\p��1���ΐ���N/Ho�vl�G��6?�*�Ci���k��0#e_�s�y7�w�Ee����]��i���4mO~fbdҌҒa}ew�&�)�^��Wo}�B�*�G=?��z�O5L����^�̪��m��ag�Du=m\%�#m0�5��V��g]ї7i��i;��ܵ�nF���_(�T����<��ҵ���m7�Э�K�l`��R�=�m���n�T�n����{�7*��PF�<��Qe��8�__�ҁ=_o�#����i�Yª��.�m�������_RU�X���{ހ	Of��t���3vK�l�w����-�h��uU�<��Q-3�jC sך//�a�G3��;_3kNa�>OE�;[����k{w�E�_��d�Y��_X��<�\���ԈKNu!q��T{�r�-���W�6+Wkۙ��e�I^3�aHY��p�*s�������oY>��4i�fu��X�^I�W�qd54� �@),'G!/�M4��CiL �01��X�S51^U�/�����KO���LF?�hGu/����O��������ܔ��>�v�������c׋��,#MA^RQ�
���{SXu�ꦧ]��pfh�ΐ�����/,�UN��
TSŃ�{��U�t[r\_9�ŏe��N��y��oglV=��㾒r�������B,;���v����N�x��Ӭɸ�o{���NF=;I27���k�yk��i�|�� m�Q;��t�F?���������ߝ�~#�?C%�ɶ�(B�ʍ��6,P���{/�u��>��4�l����^�z=��n�1��L\۟�6׀�}�Q�f]���#�i�v����	������窪����%�A�R��f�	L���1��E��J�U�<rm����t$f�ܺ���)OQ�#55M�����:g��vhg�T����ć���IE��w��8_;�:�ϴ����q@��@S��Bd,�W����]�.���H�[�I�q����R�/��{dn��Œ��BYu�aFU�}y:k�����4ܵ��2�l�h���Y�$�����wC^�ĎF���UuYA�{�~0М�@�DﬨC^�i���?�L�������fߎ=���aډ�8�
z�G�O-���1E���1c���Aǿ1��xtʰ��v$�(�u�-�L�)���� ��_u��h�I����'
..\ێ5��maƠ	�H˕�����W��+Re��B�����;�)�Y$�$|��
r�Q^n�Mv=�U�Q/:��fz����/�#�����*�[v{`:4C��t�&�'�}��=i��}d�zF�dS�6R��7�elʓ�_-0p��E;�:j��W�}t��o
#��3�Rc�A[���~�hy[R�s�+/H�?�!��?(k�VP�"�٭$��`�>U�'�k�#��(b2�����^���m���4H2�)�4�S2DsI�����9�H�>��oO�2�Y`�vrY�{��Q��i���*�t����S%}�4#����Զ�C��~eY��$�:$KI)HK�~�����N۹J� Oj����!��+m�K��N*3}��3� !)�䯳B��h<S�{�6��������Nj ����BΟJK�c:h�Q�!`�$Ff
��[Z,��o�~    IEND�B`�PK   �M�Z��?�� � /   images/935ecb41-e360-41de-b535-f88365900f7a.pngT{uXT����HJw#��.% H�t,!]�4(!
�4H#��ҒJw�4H�.����?�?~<�>�=�̙3���{��sm5bzD��TE�pY�q�+�����}�����`|���{�OM}@ �����@�H����W���f��`0!gw;O����cB�b��<6���[��O�Hl�"-j��I���_�0��p�������S�����8#v%g�Ov�M���ئŒ�\�׹�!�m���\���� �Q��	jM�3��ɞ�/���uк�����b��+�hޞ�Nܧ�򽼢��3��5$�\=Xy�{K�I��p9��定^��p���h�i�5!|m�&�bs|Ku������F�D�Wo�$�	w�H���}q-1���f{G�u9�em�HM�}v����|���N(���I�@69	�7�W�����nu���}���y�������ź��[(��wns�&�PPDD�M��M��M5���弿��_��M��F���ڛQ�mˏ҅�Y�p]mZ�wm=b��.3~�qo4��,w���jlIL�h���J�qZWLT3Y������9gv��k��ǘ��W~��l-�F)p"�C�Ƒ>m%����4�����d��%ߧ���@G�LY1)����_���r
 ��S	|;�v/�ۻ���#��Q�;�8���pm���o��	�*�\ƴ}q:��xX�Z���fE[E��_���F-�ul�C`�T�4W�0q1$��}y�J�,����X7ݟ��_	"#4��ݠ��y�M�sK-#܀;
ڥ\+$��l�ڭ��!7��4�w6p�d��VX���y��C��)��E^�=�4���
�lt��k��������׳ծ�Vv��P�������8��h�̒߬�,��G�
O�ŝ���ZW�8�H��<E(�_�a���:�c� '��vA�5��}e��P[O	�k6�
-��}%G��'�|�s��Q%�e�=|�$-3��o
èhL]�+���ė���=��C���DC��sA��WL\B��wJ�^2�jSM���$�K�:��ǳ�e3��*(��,�T I�1�e֠*�O��0�����>6�� �y�/������^D[�G����Ƥx-�6����p�*O�(���i��~�Wk=�`\�E�zЈl!R�5�y�=*:G�|Qo��� c9U�b�(�n�ѭC�Y��GΜK�ːʂn������)��d�T9fH�,:oK��<&
LF���-|w84܇ �&g��˳�骕�o�t�wӟ.m߷�n�1SH�(L�g ��v�łI*_���쎅�s����i>��XZ���'#�e]%����X�{N
��<q,U����)�P�R��FtO����v�I�.Z�&,�����v�����ۘ���Q���T���@�	�W@�u�/��w�P�J�urBp��WؗY`!�O� u�c<�$��i�&�# �c���9V� ��=�e�z�>}���2��M�tH��!JCP8>��m��"N-0_l��>bkR�,�%m��_B����S�!B�!��у4�Zo��/��`������9}.-0����c� ;) $�~�0[�ʷM$m��_l����Y:##,�� ��3���@���� ��ĀT���&�2i؅�2������T`���|�3R4Τ	�0���
Пa�~��,|�Y�y+�Nce׾�G�1��Y|�S�����ǝ��/V�=�����{`�H`����˴.��?[�T��s�W�#���X��u���4i� ##���2���o�����4�T���R�ە
B�XI������}���w�d<�Y`�G�!�ȡ�'G�*-�I��r�}sE�?j�h�/5"���ֿ��y������V�?�,���׍��4��PO��?�iX��X;��<>wP���n�0䤍�%�Ǆ���UH�X>'�$��1*�8\{�@���ӆ嶴T��u~d����N8xY�[��-��0�/�Յ�	��h.%����^�JՓ�.f*3i��p9v����"`|��������+�l*'��%_I�,P1�;�[�;a\c�mĲ7U�=���W/�
��ր���a����t:��]� ��u8V��EM�@1R�ٿ����%��x7���B}Q����6��l]ߟ�"���]'o��g�Q\�s]$�f�GD��i��gs8��s��]+��,�ؗc�z\����?dXe�#IdZ6���ob��}���c�w"��i9궒X:���7Į�Q��>�b7>����I�(SP��r*	����Ӵ]��rݮ(,��Ye�õ�o|҅c�^^+���xO����Ѩ�@
�BY4�iD뉱��ڤ��̸�i��� ����ʶvx�Y���ɷE�PNI�ο�[������MG�Q��04�BlY�������*9:�7�$��R�W�[��cP���T۴���5c�+���m��9n�:7/�A����V�z�VbA�^�ս:�Uq�`uM�09�pƼ���;3�Z|�_����/EK�g$<?<ꡥc�8R��	�JZ�cġsQ���Na�+��Q�8�K`&�'�ͽ;)s(2�`�Y�[e����oe�XҨ� a�%�oo�b��ƈj]ڸ�J�^��(x�����;���?J$���q���gML~����)��i^:�w�bAKi�\l�v4J�OLT���h���W圩���Q��s�6�S���Hp�'�����(ch}t)\4�.Hk�uc���7��f�YL�'v�z�����$����д*wݏ����\7Hw)��d�^���˭scF��j�w?X���r����N��k!8�U����$ПjT�����������^����/^<�Q��q�T�F�_W ��M@�h�vmr���ޏ�������=�,��z�%Z���a{�͑C�i[�v��ٜq�,���vȯ�s��LFMR"v�J3�EV�9�}��ܡ�d�P��'XKG��3[B&;я�#]���Ŀe2�j8�>8=-?����>��&�s�b� �N�E2�A�55�.����QD�K�Gj���i&S3#kb5�W�����c���m�Jy���ڋ~��T-� Hxmy�7D)��Ǆ+�}��+ch+���$}���3|s5Ò�9+�OtѽW%�pi/�{/7�T�����xCM�O�� �5�J ������9;�gBB���,���B���)ynM{ҡ4���Vn�y�l@Az�8С��ND��r����{a�m�څ��kI���Lp<{Ӝ��>��
8����/v���c�o1 :���K�}O�νg_�"�~u\�� �����)�0I=��h��{�qYBX9�)�����+���I9+N���ܱi|}���*Չ�^�)��RUH.:�|�^��K��K��=鵵�q���K%n��7��R n��fL�0�4.}e��" 1�F�a=u�Nbr�3i"��OA��=<��՞&�흱rO�n�)YD$��*,{Vd�v窖�Bz�F����/��R",C�g,���z� ����:����`��s\���?�������<����_��6z��%��W� 58M�y�sC
2���a�^s�F4�4����Whc���Z�9bX�8<%K���t�VV� 熒 �K��C�2�� $N陵��>��wѐ�=�H�,�2,�B98�<7���^�Q��2Щsx�9��i�]�4��+�N\� �0{\��֘�(G*t�g'm|��#�8R���~��ܐ3�>)��߯��ҹ�6��FC�.�Ǿ����9d�H�hѷd������
t�CqT<'$���W3t����x?f��G���>q+0�pL׾=y.�l�@���CS�~���N��8%�����9��(x�����"(�u�?�e��C�0ߍ?�����,�(��\�t���¸އW9�Bj�I{<ю�A">=��ؠ?4����&ar���c�ky.nlF��f�U.�҃%\�T4��,�_���mF��V�ն󷉐��a�X�����Ϭ	�F'�nc���Z�;̋�l�w�v���/�)['�m��.��+
V��� �VӶU�I�6���+��i���2�Ul�q�:��)LܬN\��x����v�KrJ�g�>�)zT֧Lk>�z�Z��x"�]�<W���M�$� �鰓�o!���tĬ��f|��ײ������Q@
��օII`�!M��otPQ���=ߘ��p�jM�|�[���e�'��8�[ߨ��=���@^)��%D����5H��)�9�I������u�+L����Ʋ�}�4�=��:oc������bX�:�]��U�k���aH�{QS	����g!�Cu}u$���r(OxN΁"�J��Ҍ�;V����ް���Œ���{�b�*x�F;� ���kH�鿮tk��#�'"s.�v�!��e�ᾥ��J�;1��"�%V��j  1�F�Jr�t
����^!�����\]�hrEj��i�m�w��W�l3���hԅ���nt���0����z�h�n�5{��;6\���lS�\=1 w{5���V�%;�:)��U�)Eٙ�+M$(��G졎Do��V���ȲD0�ڠ���oó�����'P�Bo�׮��ƀN��k֠&Wm[B�~[:��LJ��&G���kv��������A
��)��$؞7�
�-�(�2.��A�',ۤ*P�!��H��>�]abk{r�'|������˩\��R��~�
l֠,���)����C|:�4���t'�y���c�,�^�e��i�*��6絋��y�pD~WPn#����ڽ�����?��Oe=����ؠ�|:T��h��ZPu�0t����x�рo��ް��`����^	=�@:�4n�}�R�[9_�1�� g8���b�;��ͱ����j�>.�i���|;�zq���_�E_�$.m�����'
��a��\�z|a�;h���{f�zO?��!w�p8|_5ЯvO��Ү���׼���Я�ʥD�
\���+���A�VE(�$�?^,[`�;!A@-h9Mݵњ�Sx��'�-ȫ���m���(�]�S���*������x�j)�x@����E�=�13驪�Ak9��$b�]�	�l��_��A�}X�^`� ޣ�O��Z5p-�JԀE��hj�}]��Oe�^�����5q8 4��E�׫���֛n+$����T���=y�Ͷk�Y2G���u��S��?\"Q��
y�>vV(��?.���u2�јS���L�Ґ��N�uǔ&��Qѽ�J��9�	ƈ딏_�Y���p�a���{�w'�m!8��W?z�j
uv�5�� )�]ʂ��_� &#�hR�,ب[P�]�<Oɝp%
�p���c����?8�bk��S���v�B7C�S #�ў���/���nϽ��ܙ�p��?Lۧl�t}�^K�~�����9�3��rx��)����=��V���Tp�g�,f�&�F?�uS�� ��w\9�R	��AM�(�w-���+�o�,O��K0H�ro�{C����
��qX�W�{.�����H�s�}�SP�f�̹t,u�R�M�!C]�4�y��-�n�vh���"U��+WT��9w���{n�7=��`Xe�����Z��qt�.���\�*|��n�����u4�_�:za0ğ�՝�Je�&���Ԥ8���튭G�;�b���+�amt@'[S�=�~�ؑۖw��r�j�a�S���*y!Ў�b{�C}<��+�[����Ͱ>�k��e}�^�d��9�F��u̜�}��}*��[孧���)�sxv��R�J.��{<��U�3⁖If�̜��W�xqM2�Y����5)w�GRܒ� ;-��~�m�ԉ�Z�<��ax/C�g찢x�|y�wyKx/�����ׯ���0,Yݒ��M"w} `~*#tD��VYE[ � �r6.�)S�
:5`O�n�LZ��u��P�t2�EkY��iJ�l����x������h���Z�%Dq+C��w,��֎�7O�=B�3h?+RDr@-�m�C59�s�-�jBD$	*Cv|�?1#���]�Ԋٓ6����,n.����lD��`tR������h�
�740����[��z�5��J*��t=�S�1�Wٌ��[n�P��|���_Wy��:Cp���th9�����@�U��y;"K��/֡W�av�?-Y��Z��mM�p��"�`��x6���h�E��w��t��ך3t%k�jG�bA6<��@��A� YD7�^M�-Ơ�R�P&6��+��Ѭ�uB�Ѿ��W�9�WW�5�D�#����I�b}{+ZS���E�ʸ�����s�쫠_�h1���%CNg9���ؘ�i(� ��u��aۖE#3���>��������
p�V�t�����7��	������On�Q7#v�6�3�R�i�����z5��(�������e��	�d�>�I	Wo����� R�<����㾚j�x��V���!w� ]_lxT{B��V����έ����{�����W.�bf��ps���<�������~2���ߺ�m@��O��x���z�O9�w����rK�ۨҨ��<Ck�(J��;�e� #�A9\�B�� z������� ��x{�B"�9i��A�J�pe���`�ƅv���� ��6f���V��&#���d`\��oh��4��L7[��]^�^�<�.ܢ�+���~�l[��"U*ժRy��]|�!���o��G,��G�g�-�b��:��+��Ç?~�^��i��G��	Qבso�מm#�ݺ�������)�$1Ep��$tϝ[��<����6�?R��T����ZW�\1���3�J<����.QL���yպ�4Z���Ӑ;"X���TN/�٣�}J,j��twM�S�t%�5Ȼ0�ѣ;{J���	
`�z���Ӿِc�ϸ��7�ro}��
��D�F�3�"����?&� ��A����(p���y׹V���k:�SR�s����Bzh��1-�u� W!���V��DL귏�JV+�űL���[m=g1�NU���p���ϫK�B�Q;�¨���(�T��7��U�.y��f�Ba�bG��̠q+�C`�+�9��&?_��
����tU��>� ���l܄Z�[��o�z��	=�_�ic^ʕѯ���MvN�.6 ���3�8H�kU��ߣ��
	iR�H����|LO�����u�Å]��G�k�Q���@��w�dHh��d�ε*_,����6�o�K
����DJ�[Q��������V0�����PFw�/	��5:��x<��4y���z�T��P���՞�B�_ͣ%��}���n��i��͆�"*|Xm����D�
=��9���
�P_{���
=Lچ��Ʈ�U��"����IB�� ���❠Yx�0����m��@� ~��������3hܘ��}қ�0���𡍟���'i��-�))�=&Ҍ5�@Æg��&��cP�x�
��j�a���Xcy��Rf��_AJ*��r}=@8����x��`㾸9�G�����D?�ݣ�+8��a�m��E���E0ת�l�ـ[('j0��Gڜ���*�̭pJ'ȗ�3��BbD��/���~z�=���mDB����H,]K��[�d�\^��,r�	�0I$b�UV'4����Ì��7r��q�4�����c�3ǁŘBS�kw�� ���	�
�c�|K��U�ô��X�L!���+�77�;U<j�!Y;7�RIҠ���=�:c�m^��/{O��AB��o:�$yZ��\Fǳ��\')u<��.@�/���P
S��\9�c����K�깯�ڰԾmW�����o��� dcl$��HG�2�]�L�X���w�w5ߊ�L\:��|b�:�,9O.򧤨0��`?��8���S���s��!K7h@� �Ѭt���Id.�i��ÅHǴ��0���E>��y~�����j�����w��ʁ���/�ҾC�� [�JT�?;��9h��,)��v�t�W���� ��6�1%�L��>O�{�.�;ʼO"�Y�KiڧUL�w繯`�Ks�0%׃���x�ً׫�5��$���=3!L�� ����}�׾����O���>�[�g�޿t����x9����ȤgS6�/O֪G�6�����q�Z��(VQ�S�9P�jI�Nmb���h� ����4�KY["�	�|\"3j���yd'j�W�k2�����x�t6Z���n��ɺ�_~g�:N/�걭��f&@�f�;�u-q���v��^�>��Bk4�^+�0;�~��}r1�S-����BK�[�6"H��d�勡�к�ᅓ��Y�F�4��9w��ˀ��N�1 +h����8��1���p��#0�.��&��_����2�e�������Vm���Aa˟�램Y��ϛ�q达t�|�+$@�@�G���'P�N����>��5�ځf
����:��Ӿ��i�7��AO���0��x����FIF�[�l=�7��婘H����>��9��hyq֟Mt��~�t���S7E�G���8�Jns�u��!���H��͐��ӯ�W͓���i�d(��5D3w+OT��;$4E����"Ք���S�R i3rI�Ֆ yE!^Y�da���IQ�Q{�3�g�]��.�k�$;|>���,��Pǻ�#!at���2�����}�Nz�`|\��/�@-�7�& w�r�����w���_�K�Wa@67������gm�O��t	���U���F���S.p�,�����A$�'n���~0���ڵ�4��Qž��&��:< 2��
g�>�Rv���+	�����9cɔ;���m*�6��{hyN;��Z#/���H��w�S7�V�Eҍ�2�,d7%��\eT�
ha�����P���=űŇ.�+�ڸ%��-��ʪr��O֣�N�¦���/��-���|��q��P�|����׺E���6a�moSF��y�I�����nr
39����Qu=ը���,����k4��Fb�|x���Q�X��D�.G��	��������{zg_$&�ÓC�uM+�M�1759hw��[�.u���T���wF]%J���"�p�gwؓS��.,���`񚰃�'������Oo��,	o���k��t�I�ʂ���O����������IL����֦!X�7σ]�<��V�y��]�U�"�5�"���|��a����2��\5��X�����z�덁j��f@�=4'#�Fp��[�dR�{�d
xTW���,M��vŜ���Kw��I�����>]x�D��.Q(^�5v���;��ߘ?@�\�G�-c:��[Zb"a���Pjrd�z��q���v`�uBF~�i���!�ߝۀ��<���E��擎�Ykl'þ� Y��܉��6��C�ٰ����1����v�6�(��ڿ;�y@Y�f«�X�ݾ�GH5ʆ%�~K1V����lEP,�66\p�͘S��w��B�8��l-�D
�e�������R�$�O���R�r�g�޽%oo.}����j�uS��)K(��{�����%��N�6x�t~3��iA�Ϲ�#N�	)�O���/�M�rӌ��#�4��t��򃷟�l��>��WMA����gԵ1�.�6�4}Eb:}`r���x��]�jd#m���׃�P_�w
�.٭���m�F����qzzN��E���Zo�f���:r|S^:Y��o�
� K��9A�ȳh�^-}��f%�0j,O���ɧ�}k�LQ =|��Ep��h��B!oݵ>��3q��_���K <TC67���]ɒ��9�}p�i�z<�SL?N����B�׻����ꙶ��q��~�5{���r�H��q��~⌎��Ț$�@����,hфƩ�;mw���C.��*�o�4��נ\1�����P��$?R�6p�wUh���J���Q{�~�U��G�¥�Fq~�n�����9ʕa��u�Z���:a����#��G�M���m���/~������{���a�n%RH��Y�T��l�A8"�U��@�s�����Tko+<�W��)��|�+!��r�ɖd�*V��K;e[+
E}W�?�:n�7Sas��LS���F��YkP����.��z��џ�v	q�ԡEo���0�;�"�j���!�p���D>R�)dI�x'��R8�W-�V��
�x[ݚ@u���d��
�nZN�q<BA���G���^�i�]~H��㊶�q�XIDǏ���ꌊ����9�5��}WIa�6a���zE�[ZZ�C�_j������F\O�Oϥ�	[�<_���@:Y�d�#Vh�H�H�,$�+uo�>�;�4��씔��5l�I=�j۟�Q�!h5v�Y&k��ݬ�^����We��KD�(��="�@7�~b��rF�ܤfE��a;<�>�v����y��ܯ��`��R���JR:�c7%">j�����2@
p�7�w��s7��a/��0����0�UNO���F*o�Ӱj�>���j�z�5�����#
�z�	�i0�3�`��z���*nq�$K%�l'2}��������SW5aw��QM-vS4���k�/�@u�����oB�f�&39*�[IV�w7�Ĕn��X���yy`�k�&�)< Xt�/�ۼս$g��7��d�M ��齈��+R
*I���m-ӹ�oW|��s�H1=3�>y����Y5����_�����EgK�/L%��Cy���a���go��Z��xP�\�ړ^ۨ����
M��I��Z5��v�7R�q4�1�̉��Oŋ˙���g��L��qW��;���r��8�٩p��@�0��S=����B<���{��j��W����[��`\t�cU��Y=v�z�J��U�ҩ� �l�9���������7։�j��'xX�� Z����h�x�A���)R0�h�y���q�k"����<��Ǝgw�1�'Sw,8��0 �X�QNp�'�e���yu�rm=��sl�$�F���ڑO�-p�T��m {�={������Qؒ��N�~�Z\Y��-��ݭ	';�]|
��[��<������ 5��!ƍ��+�]#��>o����y%���B��Lv�I�`��\�[֦�a_@�"00nB���-[C��5`A��e4����j*�|4�ҁ55���W?��X�[�nVN�T"�BzP�����'%݅^/��h5v�ު��0~��i}���h�� ��#���5RLZ�fs)�����H96`����c��=Zt�\}Jw�� ���~�6�ȏ�\��v����yHp wqußn�k����]��3G����n
��|�D�]>�#+���=�5=��38Y��K]2����f��
bcj�Щ��ox���w�ԙ���O���8����M�;��4#�g�
k~;Xg��<�����ӓ��, ��l������%��q�ykJeؿ�{L&"M���{��l��ɍ5F���]_�P�J�$ױ�]|�Q�a؂	��BD$m�9l�m1�n�^l�@B��Oҩ�{ޱp]!?Kؚ�쇐r�^��ӓ�X�����]T5>q��� ���y��ǵ����L��s��s�oZ���r��gb�������w��k���G������[C�'�Ȓ����N��9�na�CV:�b�WIrb����� +둄>�UP*�����[�Ѵ���&]y�.5>��C?y�Έ4{Suf���Nuy�!�9;/S���pP����T7J�A�����7qqG��ZDR'���!��&�h[[I�����,O%x\��{~(J���� �5t;
����|8��r����l�x�-5�,θ/�UX�~2�O�U �z�Q�����'��y$�X����<K���X(W��)4b |2�������\�� #�<-(#~�[u�|�jn�f^�X����*ܱ�mw�����-�g@*�(�S��{q�N�}�l�7�H[��;{Ax;B�`x�ӷj����D��,S�4�L���Z0�^�Z�����Ԗ��>U��1߮�Kr��DT�:�3)c�~�2��ͬ_���}�Cu߂�v����$�1���|Zz��/ �.�ȫ�E�	�87����r��. ���� ����=�P�������UX�P��o\�bN� �r�̞9.i�+4O�/�
 �EWx����z��B@� �>��]�@�t3hZu�*���Wa��Gѻ���YY��~9���F3��xo� V<�(r �7��g��Q�,�8����y�=c�7�}�ޏU�z��w3��m�Zk\D�j=r@�����h+x�-���Mf����7�v	�D(�Ry#e�>���WFj�%{qS>%G��)�)�wh�׶����|)=�	��}�$$L�*���M���<l��,I��]�B������Q�`�k\�fC�Nc��tD��w�y�#a��b�B�'�e��	��X���'�k'��ჩ�hɆdIowWi*��2;x|��
��ѭ�d]?���'0�Q���O�ܠz��V4�#��|�P�/�\��ސ���ߕ�P�S�`]P4m&{,H��ku5]Ӗ�^�uXbD�"�v��������g˱���4���c��\�s"�G�lU}l��h7�5���y+{����(&F��&Df��?�Y£�v�-�cTa���sc�2s$���7�&�@$C�����wQʫ�ni;�u�R������Q��z�k�9/8�yr2�sh�a��� {�?��@V#��z��N��ȫ�&v�������&' �J����} �} ^isLV���y,���	<e��UzN�S�*��f5��=�L�-;��mMf:�&��,�ؔ�s��m81�mn��k�'-�N6sWi�t�D�� 9���v����3l(���F?S�}�(�Ck�I��
��P4@�th)8OJBoa����I5�*W�v���F)�t�1#�[h��p�	�P�)�s6�Uл$�0�8�~�^�LuU(;yr�]�
'+��
���Z�"P�y� b��܊_ڀ����8��?fCgNw�_����-%�+{�_���+�\׉����#{f��M� �L����
��b�j[A�來�ş�qHχ�V����A½�9���Q[�lP���Y��=}�lQ��^ǻ����1�`$U�$�����MW��uC��㐎L@/LrB=C�DT���P�*ܔh'���Ϭ�18�2@��+����h>�Z��GY��Ű���M��x.e,pQ�������H�?�~����}�;\f���a�|�3	=�iLv=e���gXp�8��V��C���$�ِ��(&C��!.�O����{��w͉�n�y1Ij���u�z�u�<3��$\�o�Y�@ӝ��6�j���auhY�ғfMP� �M�<���GCK�yMˋ��Z��ŚL(	E{|�BO�➌Ɉ�ԿR��k��m�|g3�5�I.���uf'ֺ\��h��͑����u�Ʀ����o�4�e�}â�Z���ϥ}F�wW=f �7�y�u�[��b�t��f�ۻ�J�@��S��=_C��j����
�����t��\���F�x���<@��
:O�J3H���׃��i;��M�ު�e0_������{��m��{z�W`|��qu^�����c?�Y
���X��k|�����/^�0�OOex.��h%ԏ&�Rv�H��M�D�P,!�y��!q~��3B� ���3���ϰP�7(s!MN���~�Oȯ�p�I��ep4\��
K�о�_��3ɸ�W4k,�Zm%î4�{h�z�Y���"1�����'�������s�j'#�����,"�0Q}�fW#�M�1���U 9'�E�!��A��m%#�}�M|N��D��
}h��ي�{�z{�߰�}_����N:��5����D��YЩ��Wk|uVհ��@�E����4���5=$�|~�zЅ�ݭ4+;�C����cM�m���h��a2�q��;.0V�iI)X���	N5�x]�����:e�S��a6�R����/엞��ϖ��M.ؘR8B���sT�b���I�<#����'�6�eT����#ۤ����:����>�s_�8/HڔB�цaǯ���������ҐM|�⩄7$_{�t�Im��_k��.�Y��M�Rʮ3N���/����-��_�����3�����rE��	�7��*�vj����1h��].hdN~D>v�3q�¾���}���N���X7]�wZ�1[�bG�;Dk��-�˱0��r7�i򏑣��v̞@n�ѱ.i���h8pذ�x��$3�8���o@��H�14J�}'_g,W*_ϻ��-`�~�c��k��1����:�	1�z
� *P�x�ٷz,'9T�謏Q+	T�}��C�U�&�[�JQ2��:��\���Uwu\r� �K{zp#����+	>5g���J̓��g�kj�ǭ])��2r:�u��:�[��4��BO> �ES�1h[�ҕ��ۻ����2���� 2Uش7['�$�u�i��B�����ѵ?�7.ɍ����\Գ�anE��M����2*b�������Ì�<�jO��3L���z������8ZsP
�[<6h0��4�M��"�sSr8�?9!m%Ul�d��`b�/a�;۹�G�֩��SbF��x�w���0cŤ�u\*�"[���=�j
���Z�@O $�s�޼�*!����.�Ox"��R!�1bT@��G�ˍ��`9�	���>�F�=�+zP��m�ɢ���z-!RY��:O�uaeQ��8���a~�׆�>�F  �z����=�o }�5���)�A���^���|����N��{�]1��|	�=eI�a��f���ѹ@M���_�ԃE���^�)n�'_Ln{I^넁@��G(=�1V��`NzI��)�)]s�_�yIH>Y��=�P��t&��| ɦ�e0彗��/�Od��AF�n;
��T�+-ޭF,���x�g|�q%� c�fJ��q���n	䄂Ll�lA�J��	�<i�"(�A���.O�AD`��Lٮz{z�z���D�bh�&,c� ,��~��Sh|b��9i��� Um��N5̭w�:>�Β�2��-�ȯ����Y��j��+'�~&��}����	d�\� Lk����6�PW�(�m���>��,�[Y���Z��_��l>�#n_ Y�pJ? `���1Q5��!��q�����i��9U���o�|��U_o�WÝ�����z�"&��*�pcZ5�ъ\ 3���������t�0��og� ��~;T�����e���{d�^��	�Ԋ� 4���� U�����,����#�+�1�bR���Q�@����#4(%8q<�@0#�Y���`�"���ɖ�������u����r��7s��ܠ��6*E؍���Ta4�y�fW`/�3��oҾ�W��a�M��i�~�y�Ԡ�ˉ��!\��-.Y�����R)[����^�&Kr�Y�\ NX��QϏ�i��[P�="�{ir�L �����g�l�2��~�>j3���2���<���y��C`#��ϸ�B�v~�'��h�|�1� Q���M.'�ex��Bp*ϬW��a�� ���ڹ�]O_{���]7�S?�
D�l��<ɨ�������P\�|g�
[�1g���7Q�,���>E���-{�V�Fi0΢�αe�����|$'i���;>Q�M� ��D=����(�(��?;I�F�U��2j~�z���5m�w%¯��ŖS���Vy�c��J�+�k-���=pҠ�x���1I,6b���=�x(��� �-�:[(8�%���������D��A��N�+6߁2�d���I��ˈ���V�����i�"-�u���-Y_�_$��]�S=��bH�?|�k�s��]�������iG�����W~K ��G��GZ�-+���d:��s�ˣk��Ǳ)96�ƞ��_/C���	��E>޷A#�X��]�s�P!��9��&���D�e{Ax�0]8H�_�1�q��lH,��9AN��3�?$�~��vg�5D_��� I�����!�߮�(���\�I4�ZB�NV��7>f�������W*v�Xٓ<���hڑ8��x�z"avS� f�IFѧ��[�01�����;%�`O�g1aF���W��9 l>֓.}����kT쁼6`�M"R�# 4O�W~	�����\ �ӵѸ�����g�̅��fxb�!�����?O�����B ���]蓥e���g`��j+$�U��5�q���/X��y>Q�|��{/�!���類�HE#h>�J�ɘ��>�3��T��+����X��gґ}=�������Ҹ˸�|��_Vk'WL��y�:�:PJ��"��gf+A�M6�c]�3>�⊰ٚ�UaxGb�z��9oJ'io|�N�?[�!qS\��w��`1�|���6Au�����}�4e6Ҁ�RdQ����D�O��ڸ�,���e���������+B�C��m���7#��eŁ����\�ٔ�������C<�t�QX����x�H"�oPh��:���m�Mȋ�B�M��_����Z4�c��r@��ȸ�����ی��T��B>��`�1NϨf�������(vK��g������:��>��Hz�[���Fgܬ��h�u�G��,�2B4�����o �j�|��!��u�ԎTu�	�Eݔ�6�()��g},�y*�"����k����
���}�E��Z&"�Di㯟�2��X)�"�����*���J)�n�Aiġ�CJ)���D`�n	���A:��n��;��{�}���ϜYg�^���xUD�%�	_wfb��'����Õ��4V,�4��h���7_�v&�G+&d�3"�t�tv~�0�j.'L��Fj���@'P*�*X�I^�������p�`�˃�	8���]朆K%�W��3՞6.� @2V����+�0��� =y"b��D�Z5 O,"��\�D���y��]L�D�����`��8 �d>%���}M���mb�`��*�~x��.K�M�7:�@��FQ�m���h�}���J��
�����`����AoÑ��Ĝ�� Pv"������+�0�YB����jM�K������<^����Gc�F�M���OƯ<\oH��O��=D�V���z�1 0��k��	4������W�3��F��][AD��(�@���J�՘�0Bs�
��o/��H
@�`~S�W�U�����aX�D��tSAQ�10�l)�4!�_L`I~P����WlT4��z��~3U�Ȗ�֌X�n��)E����dF<�?����GT7'Q�We����!]��7�.\���j�+U�[%�����)��\0`��[B���̎�-�Z�~�)�)�`u��Kr͖4�%�|CFNm�kP����A�Z�~߼��zj_�O�P>�����w��CO(bM}B39��P����@W���A�\��C�Y�1^�cv��!o^r��eY�䊧�u��h9qx�k׳�?�y����6�-6c'��Q㹶�s.0oZ��Q���ԬI�c�	���~�-b�:�֔�|m���X�v�����?�?뙭�M�ao�Q˴@gX%R��I-�+A�{��N�2���2�	'�ÏR𩓧9�=C/���>������f���`����/l}��
�[���2\�M	��t۪/�}��ct�w��m�����7�Е�����q?��Nl�&C@������QQ�m�9r�=4.Q��LS�Z��"(����Y�A$�X�n,`b`(���zR�;Ve�$�Ez���/���k�P,{��Y�HoY��\���/aJ���l
龕D�%Y��4�߽;��l�#��?7
�ُ�6�$�}'� PI�Hm[�α�t�}#��S�y7]Fo!Z��u���HL)Cm�\T~ɴ 3�[0�i��(t/.����lj�8�e
�Z���)��>)E��q�J�i�i�F"��8>r�ح��gׅߞN̦���s'���M6�8��Wr�+�oݤ3#�[ޅr/Hd��sg�f4�Vf�%�R(��*J#<��O� ��WGB��Oo�i[{rW���8��+n&eh�ymh�؄�1e���+sY�d���rsL�-K����zue�A��c5�|�-�5��5�_t���70�
�~M׏��D�4[����)��1�hyR�p�&��|��Jw��S�~��P(��� �Y���B7A�P�f**�F�,��i�Yl��{���2������|��,J�g����h�.��>���:oqt7ո��wm�x�틱�&����fE⬂�������W�W$��n.F.s��E�bt�j����RrRRRR��i�^�0}���.��l���N��y���������y��!Kb��.Ih��Vk!�tP���Գh�W��B(\	��r���ە�w��R:%��T��S�d�M��W���BwT$w�]�%)྘�7��pg�%���Hu$��!ue�ȈY4�oz؟+�ҡC/t��v�żT`���?G��Hmp�h��E�{e8�,e��������gg�(�9��!��|��ScB|������1�ڎG��պ�]T��pˀ�^q&�o�&ٸO՞EX!��'�����/���dF�XH��J��>2�C=>厹�Ԕ��?�u �A^�wx��S�����?��*Q�Q�\zv�C�&�sP�n���.��;,�];,���n����$=7�>ǹ?3p����U'4�޿�2�;I��+��1�s�S)U8+qo0D$�Q� �0:�P)M�KL�Č��/)[��6q�~��c��а%/�W_�P���gC5J���f� ����`����K#�ޏ�%��9Ev?E0Xp˂�I��V�+.�c#�#�n�9B��_7�e@v��x	����^��,�7��T?ڗhvy�AX0yw��WCS1��>�3��ՙ��ۨȌL~��}	�UQ89�A `�xH`D��G��K�x�ф�Bh�$?�M���>����P�#w�=���f��<5y�c8�{���`_�8�z}��֧��c��6���;?e(�����쒷�]&O��GJ�31~+�o�܁�Wm<�rf�[o5��]wi���kȠ�M�P}�L�����B֜���W��ë����]�w����̑���-��L���m��Ldmٕ7�L���z�*Qc(n�3��m����!�� H�,��Q��`��za�lT���Ety��֏�f�٫��P���E�~$�ӹ'U��j�<c�7Q͜����s3]Z�0{<5�a�緂!ZA�!&k�9j�R\΄ʾӑ��q
��8���;|��-��;l�hB�EjP%��1������\��[*������n������Ak�d�������+s��CA�&�[��ZZ��P4�c�-.�?�Z�,�>�hu��O�ڴI���m�(�6����|��޻����)�yoR�����%sc��J?zg?�y�f� �z� �E,���b�2�a�+��Q\i������kL�`�di�'[�>�31�y�0!�Q<��Fo÷����q�ʚ��g�"o��u��Mg�4��酥´��zU�N���D������aZ�jv(,���~�������j�~���颵��!���S�]�R��&��N~=�6��vۂh��l�2�
`\�NFrd�9���Y!y�C�t�3��8\]ߺcj��Y!+��J9I.a
���e���v}���+68�4|S����M�I��ck�hPr�*�w���V��A�\�a�Z��Ѽ^��d�w�,1s�C�ץ�V�|�9|�"5K���9ˌ�^dy7����Zx}%������9C�6$!��+�%�փ��F��\�,�������pY�Utf���������0,�7���o{��3�*s�U8LI��I��͟�W9��KZ��Τx�>�;\2�8[����Ѻ�ߚ �[I}�M�,fq��]JB��9���re����c�ϑ;ݝ>5����T�Hk�x'Kbc�U�yeX��nʓ`�\�U.L5�)�jE��#�o5e�ǜ��m띦/% �/&�k��nq�R�˙�6�%����I:�@�S�P͛/��mz}�4ȯK��
�Z�mcB���� �ɪ�F�l���UM7��9��9��jO��|�pS����]+yG���,�CL�`��Ȑ��$���Z�}���Fy+�U.j~(x�߰�|2�c�i0���Z)��nč�l�v�ܓ��ByWwZ���+Cf$�[�����.�_F#��t��l[�$�kO�o[B�1v,ǖK����?m<WQ�"s�&�~���m��;�_�K�m�(V�Zia���j^�]N=Kvu)l�ő�]^�)类�Y��љu��574�,�}q��J����v��i�R�����mI��m����>o�5�2W@]l ��_L4Ṡk.�h�#�Y~�R��/c���O�\���|1F-��n~<D���fۊ0	�(")2��}�[w�mt����[T �p�Ie۝��u�39����$B
��+��xYY[_w�T\9���}��iW�"�Л�ڠ�cv}��0u��ml7�t���h�����	_L�I4�b#��"q��
>�+zւ�VG�a�%eAJ��J�#�;~O[���ؐ#�pY��o�����C)�L�6D�s ��if�#�&qI�D��9�_tf�=/�~2��N��bƲF�ܝ�Ֆ)��.pm�!0��)�'�8ۊ�ͱLP߳�zw��F�/�]̸c?���R,Qoy�m>Y��)$:��a��88}͚�6�G�H��G%Z�OM�h��~E6��bf�*N+��k3�U�礙��ߚ���Ơ��Fi��w���'��B�&�ƌ��T"I�~��X_��a|�����`,���i���|[�@�֤��2�Y\b2&�( 1��l/�_ݎ�&��Ӣ;\�G�f��Ԧw1f��e�ya�ܼ�ޯ�������?�a���`�vB�2�������(dr��;�D���ń���8���bMe@��щ�q�.,��,I�uU<l>5�s��7X�����9����p�E.�JYȐT`P�O|�@������*h�Bx�͂ (��u��j5�#����v�qY��DRʪ#�/����P�dA��%����lzP��/1u��Wm�5q~���Z�gfͥ\a�}A�L��<���q�^O��) �7�� ���M<�\�p6"(ۊ?�0݌e�J�JS��:?x4D�8D�w�w7x��c4=%N�������� �1�zu1��-m[�
,�^��1�_.��aV���.��<�-=+��׀�e���(�Q՛��,���ŐG�C�����"'-Bc����N���5�V� |)E��IwOWmi�7�(��,���Q4Z�PyC�˂�5���ic������6�4��%�r�����}=�򸑄�k_��0�x�3)�A��礷s���/�C�����ʋ�ޏ�ۈ�v�C��o{�@�����|��j2'v�m�`����S!b2����k�IU�wi8�.^54��z���6K���T�jo�,�qttN]_9�7Qi��?�u��ݤ�}OM�0�&v�iM�Dҋe�|*�y���;�:,���C�$muDD\'h�v��ՅK:M^���ml�f��w��I{������[Ϸ�w��ᥜ�j`i���%�ڏx�Kl��N��<l�z#Q�A]Se�r��~Qva��&���I[��<4���kq��M�6D���VJU�U�ʷ��vW2���_�3�]W��`0ڢ�	�!��BH`�K4)-�[o�v8ϯy	�"v-X�N��`Z�0s��^6�r�f�YUh�\�8�M��+iع+��p��]�x[���ݬ�:L���!WL���[��4~�(�3I`M�$�3�N0\Ы��ژ6>}a���ڲ��O���.���0�L����ݘe`�},��ڏ�D��P����� Ll_�Yy�X���5�z��a��j�K�'�ω7t���xm[��k��I�=��^'b�'8�� �+���b�<��I�6��e-S���4-K�3��~s泴�ͭB�{��"zW��&�}ϗѩhS�o,[�H"�fCSvl���$�� ��,�A�X�8���l�xذ��y?m����BV�c�uY9�n�B�@�̡Ek�;�5ӗ��#"iy��/X�Z�@��m�O;��2@�`�0�/ƙg�]vO�>�V>�S'i���[�Ek��-)���g���|#�"/����V-��馀�wHz��((�u�y�	9*0[�IJi���bu���$G�	�F��l?1�A�bg۩����\���6��w�5q��zb2ᘧZi6�J瓉>�'c����`L���mA�[ۘq�<ȍ�@�X�;��M��t8<z������4��� "�>�WnC�y���Խ\�Sh7�6��!/��t�_r�\@��@h�� \[��/wd�g���;	��.n�b�jt�����xj��G9�&%'tҹ"(��̬��G���u[��8�s�^�B��I�1�ɤ}�FY4��!���y(|�Q�vj����ҧy�+w���Q�G�~�rr�oȷ+O���n��������]5S��P�
��<���O����d!�<�Bb�3m8󒕘�ƺq��&Z �2��2G�q=\X���6F��i����;�p$�: �
�86��C����	��v�Qyj8%�b0 ������At�.qB�<�U�`>U���ܴ:}L#|R�%NVD+:�����y�L~U[9���?�L�5Xb�IÈ��$��z(~�9��d�^�Q���	[7�EW�̿1x�����?�F%wurt�EK�b�X��W��>�t�YK�o��J&T��6���A��7�	I�&mވ)�4#i��c�Aٳ�o�A�.u�;'�� � _�Mδ�/���>#�������ޗJA��'�0�˶7|�WI�$�z��Ѧ���9M��
ߴ)��[��$�B��b�td�{?�_P�����|�46b�7jOnRW\1�7:�����ą�"��$����"ԇU2Z03O2�Ӫ?�ۉr����>93���͛]0%K��LZ���D��[Us�]�����d�S�$%�è���3��
�}pછ�]�.J��0���!��`�g��p-��t.b���"G� 0�u�v �Y��0�z:������1�Č���B�Z����_��]A��>��9-ڷ'������*aXV���WI��J���2I��{��0�q�?�J���&�k~���c	ȸ[
M���}��u~\p��M̠�^5ۯi���eJ ]O9��l�A[�}Z���]��:�[�I/	��n���)I�a����³��b����6����v���ϣo,�N-O|�}�>"�������4�\#����� �]�q�	��F8`s�����0�o����N���H��X�͍nnlֶ�r�b�ȍrvZi���x���W��Mq���+�T=��>����]����鉋G�0��ڤ>|^�?v� ���%cs�2!�zO��JW=1��?��a������I-��t^"!����+s�'C��]ө q��<��*�:�^n��Y�������պ+9#f�2�iP���^)h�3~!�n�y"z�y0��|῿�ܓ�9Cqhݽ]�J�h�l��~����k � ���$�%�]2k��)b�h�5��pI�] U���q/؈%a��ay.�Ϋ�!+Y�X;{��J`�oцW�u�vt��6�Ԫ�H0���=r�m1���ޙ�';L�Ӣ@�:)U0a��m�)C�D*������00Z��u[%��/TբKcg�R�/�럑����T�~��v�������:��J���=�zPF%ԁ�&�QW4���\]s��?`xy�Q�>zbW��ӵF�g=8��A��������]�|�%sһ=O�&,
�R}�No���2���8XYʧ��!�Rv������u�g;y�,�����{,ŖOy����h��y45����������RN�H�{��ɥѤje8���)6l��BU�k�γ�^���E��x�� ߟZ��(��2�(]�?4͢-�����1r(.���YWv}�k�SɡP=������������5��	"#R2�S'�^�h�9���e�3N>��˿ch+�{v��3�fpiI@��'}#5iuSm����tִ��OĮa�*���o����� #p�`�m)¸� c�`��C���n�Eu�0�T������Z	���:C�4b�nϒ7��)�� �<�}X\^�
�\��q:�..�����Ǫ���?p��~_��P&N��&�j�R֓ӷe�a�������p�3p����.��I�Ƿ�í�8�7[�}G�=����z���8k�M�[����r��`cw��ih!��Bɵ�s�+�QU�݃����z�/?-�W=��
Q�x�Wǜߖ0\s��_m���r,�5��O��9��S��A#����{�)�'���)��{L���`������e�����pl���2����뇗v�,�!��?�� �#*�Kz(AAp\�;��|��a^�G)K�;�+�P�Cvmu5��;B\:�i�'�2Qs�џ�q �V� ��� Š?��<��<�s�j(��q�$��e�x�+ЖM7���i���J�"]>M�k�~�ܡa(��m��x��^ս�E�'dw��+��Q��m��|�>k��n+�i����R�����t�/����
��O���lI���������x�fǥf�(�9X���F���f��6�MI]A�An&�?!���,&Ӌ�iUDjڋ�Bm�c)~� �9&��1 �N��7гb�/��
欣�C�E}fag�Z7�n9us(sfy�Q�ᯌY��%@[��F�o
��YZ���U[+,Rj5�6�(Dw�Z�qz
��08�C��̾Y�����T	�H1�A���)1I� l��:N8�70w��M�dBH��M$-��X���#���P�׫������U�C8Y�=6I����'����]ߔ�
���۲�%߾]��%BŦŵ�ڙ��������,�A��ed���-���oNz1��
(Y��1�7d/{qXIy��a��¢mLe�6������Rb�O���x'�_><���LuM�1�_�B�3�>�ϐ�P}/�m�[��?�zg[<�2�����w�
R�?�f�_Iw�5,��q`%��_=��LBab�H,�E/�K�d�^�D��<��}>HF!��!�7�C�ϐ��_P��F'�!�덧��O�,q����6��<��^.3����JL�� *[�%d�S�^� �u� C0��tq�}ʻ~�����5|P� �k@G���WC��P�EO��A�Qֺ��eԵ�(��	�b�����TU$'���nz�$K_�>g��A�G>��
v[�k�H���oK�E�]�rf��oĺ�wN����� 2�ZZ����xǦ����U,&E:�7�l�2WC�[y�}`Hp��$���A P�љc�2}����0ݔY��c٤�����_�$�ۭ�U��>��TqA�ޏ?�	u�(J�ƽ���Խ]���Xl�g�(�{�+Uv�bwL�s�Ga����@�J��<�2�F��3�����0~�T� Ͽ|><W*/R+&j8����YH�%����\h`����[�P�����*��i�[wh�3�/�}�l�k7F�����;��C٧H�k$�ӬhJ_	�[�)��4F��N����z�w��4
��1�*�jxd�J	�?$�V��ǶkX�S����A�&˰��J*�]�� J>�O�"��Um��W�9óE����׈��V|��vuKX:�,����BC�Ǌ���%#�m�b.����ُ�FĿ+]�;��c۴B��%:��5(��w\�B����jӒ)�*TE����S��iX8�P�)���YBHH�''ð^(�񢸋��Uo��9�ӝ�r�u
�E����+�po�z����-b.�ޣ�+�������E�h�ۃŀ���Ƥ�4���:����5H=3�s���&ĺq��ރ�����(h{�2;Wv
�-%a�Y9�#�0*~��tM7w0����XZrzm��a�Y��ڌ�|�,jSi&�l���K�\b�;\1W|j?��f��a�AB�B�h�z�/�5�u♋�w.a�M֪q�
Š3׽�F[72�M*��}'C����"�x1��H2��Oo�5Z^���3�A��v{�O,���)H
�J@�)�@<
nb�����Z>���Z�)�ġ�����3�y!C���~9�Mg�n�t?\2���ǖj�/��٠ߧR5������A��a�'\O1����"Gj[ҿ���z�j�{�W�(x���թ��Dh䨞{]M�������//E����t�F��÷�@���.r��Ś@��R�u��K��1'RkΫ��s"�5k���LL����<Õ4�W2���P���\5Ȭ�� ��wŐ������<]�CW�%#:J�<�0p��etB�xl��q�:tE+ۋG�
�QSq�l_�I����zS�V:�G�n�>���ځ[vT|��)گ�JW��0qG��.h�.�d٘H��^���#D��gaN6�-�*��i׈�4Ȓę�*��*&pj!�41	��D �s,3�N�(]X!Z����aX�2&N����
��.E�n9�dR0�'�}�k R?WD�3R�;z�xz}�X�C:�^_�j �7���	c��7�aO6�(��d M�x������ϊo*������/��`��ȴŀK����Ȱ.�J��]}�vT�=�H%�=��{6l��9׻Уv��+�J�m�A�T6]�-w&�ҋm-R9���n��d��b@��Q�#�Nak�m�6O7簱`���B�'ǃĳc?ӄ��	�@��)�<m���L�I��g�c��� ��-��LF)�h-ɞ��v�}4��М�~=�i[ ��-��j��jh^À���E��TR}�ݬIfl��ǀm�n�`q���ۺ}��Վ�[����(�øyz�;����đДx�n�8��~(l馳֧�!���چ��n�'���/�.�j�
x�۫bIc�7ݰ�i|[*��ō9n �����}�����#�~q�"�p\;�o`�&�`�!�q�0�ݐ��<��;�f����/�q9��^�{�'ߙ^:�sc
�/�y%T�s$�
s�YG����Q0���+j��(Z�I��@�BY��)�y�D�uU.ڭFO "��g�����34�y�qש��6���h��i�s�ܘ�9e�n�zKſV�0F���.��<`[�2 ���mR�3ymE���WEɠ�-7��ս�/�d>^P�Ԓ�'��?��T���z���j�Bh��{���i⟄��I����3<!���{S����|H��D��WqZ�Ru���ݎdX�s�ͬ����8"������r��N#>r\�k 26�JD���x1,0�ys�H	�xڑ���Ŕ�8�=^QY��Wt�>�ݟ��4�]F0h���)l����ã���P��0�.iI%��̎��\�E�d��c��t%G	($�،@� ���5-lx�$�d���DG8]��������UU�܋�Q��&����!K�/���]�a�"���a7��#â Zd-pmfd����^�s�2���!%����u8C�>~��F���!�k��^��z��G��p�{K�H����;�:�g%���J�F����9
B���O��#�;y�,�[u�
d`I����N�<����e�\]�8\���3N���u�-�]��U#�2�i�UJ�: U��ͳ�<��;ףw4*Ɯ�wlb��~�X�����g�C�gg��抛�m%+�<N��o-�Z��-�8+!k�'O�d{@�3�w���u0���7���ԝ�?�Ń.x|BK�"?��b]i!_���J]�o�`�,wt��A�6����a������oԵ����ƈ_b}� �6y�?f.��ըSG��C�Vq�ל���'�)���Gl����m�g��Z�\��ウ�[܆w�,�[��[M�5�w-�Ǫ�� ��2T�K�.�)l����\e$�q^~B>W���3V��]�LN@)D@����dz94��H݃Y��#]�k<��ނ�v	�3�����G�SE���_�7�rZ+�<-���Iv֧����Q^����L%�꿚�ȿ��hI �:	�^��I�~Jjg�B+%�Ew��`��|�
l΃�`�.��|���%y8eb�̾�!V��Y4o�ۗ�2n�
d �O��k9���!�⾄�U�%��]M'g�iV���w�D��7㐌�s���'����v
�;Mc.R�讁w�=>�����+$2���'�a��W��c���ټ��!"�c���2��C�E#�♢�rf�ټ^��>���	�=]q�yVbٯ9�x�v��v����Q��<@̔X��ʾKɫ��;z���?E[qD�� ��1��t^$�P���}��NZ#��f-8�q@9�`s�].����钷O����`����\ѳח�����s�&��|�g�,��_��hV1���y�mԬyq��S��%0���(:/���ۑ�g���Y����p	�[7�M�9ۮ�7��jと��f� ��X@�Ť0v���w��,c` AN��-�d�縵*[�q$%�liV�U�;�k�rm7�{�7��	���7�#S{m������Mɝ1L;F��蔌9��#�"�ɚWf_�bS�'>g@�,��,x@���;e�Q~�X4w�
�ɀY�~�h �p����4Ӹ:=��O6n�سe�������0���jP2��GtU����|��\���)pb���P{�y��Ҟ-r�L�JrYٓ�[�LQ�!�(�Ԏܼ'�o�+��V��sٚ{�o�?�/��U��o9r�'e�������@�^8����z&���0J��;�.ӹ�K¨6Q�&3�j1����Uwd���HA�"mK�>�d��?ɱ"Z���!�D�#�S�
D��[��˴2�UI�T�Ý�w���C��RD"Ӏ����00<>�?��N����L����#�h$S��"4����&/-	5c�\i���KJ-[W�����胗[�4�^��d��S��Ap��5��C�d��D�-���)B(O;EnE%�WW�M镉oo���)�dE� �̫��6��e��Â�Y�8��ɐ�����1�)�9|�$���D�{}�|�Zy'C*�-��nB`���	�'�Jq�M�<�f��
ϘfB�3�.�z�S�K�w˗��`��`/�}U�������5]ګ�׀c �E�$�l��`�Nq2n�Z���Q�{{�]���r���T#�d�X�Ю���M���+�n���6חS:���?S�Y�U�ɲ����:���������$� ���t�i����d��-%ao���֗���ќ'���D��=WS����(jY<cہR���B���x[���3�!�#��4�)�Q�������X)j�P��2�^�x�5��1�\��j�~dt.�A�*��1���`���rE#��ԞgF��?m�	��敖�4�q3Am��q���x�j�<J�m��	�v/|�3��G�\�򗞗?�W��h����:ئ��}h;?���6EV�9U.xj(�1�4|oA�������ċ�Ȉ.90�Ͻ��������c���J��տ[�{��o��{��/:7`���4�2R��8�����
�c��U�����L�%oX�8��6~�f��l����da��/s?��L��]��� �Vgб�]�LE��2��D�S$G�3`"t�5��ց˭�_|��^�W TT�GVh�~@q��Ȼ��C�����4�c���'�D=���w>�/:x��ֆ�Ӌs<:d9$`�3�8D�kP�:	��0I��N�?��#w�\��ɋxT6�7[תA6�u�(��í9ͧ�B��#�����
�����]1,ו�`˒Z�gWTܷ׊=}O���N�g`�n�6~�A4$0[�i0�O4}��t^p_�A��H�qO��ǩ�q��{�j$�!�v���ӝ�RR�@��ec�fT��uE�X������!)-���gb.��E\�ݞ/����*��/g���ц�o��Z�v)E<u�Ѝ&�:	��h�Q��|���ì%�{OE�%�}�X>�e�'�[$��A�U�P�/8��+_���Ì�Y�q��1O���f��sl��7CRhz�@��U���B1������<A�]��͖�0A����{\Tl��D�2��2}βWJe������i5�n�o;ӵoj;�ϻ��Tvh8�շ��t�|�>�-�!��u�z��<;��o�3�A,�c�T�{b-�FI��}��7���K~��w�
��-aTm-Ʋ
���K�������MKΖ�,Y,Fz��R[]��<�(�V�×vy�M�88R�rxZ�qH����M�aN����4��+��VE�ĭu�Z�&Т����s�R�O�vC������wJ���qEt��Fi[6.*M�O�ɞ>��j�yZ�ɢq�N��@M3��1��S��g83ւ+:(��5vtP�kk;ι��^R�}�\�B�پ���E&�H�n?�0=5�B�'f@���?���� �B@��h�U��䀤�/ѥ:�;\)��ZU��п"2rʬcu������]Az�4	"���H~��oL���}�?<���_���>���k�aI��{��c�-F�&$ZV��&�#V�kF�8��.����U>���d̞
�"�L��҇�^d��t�3T*^O��'Y`�)��	�����i��1@K��vO�y���� ����,D��	�������6�Z���s� )����U2.̐U$z�}�HHW�����A��<"�%^t:	5<��x�.l�=q�������!� &4q�~4�vK$تn; Yܿ'9z�+0�視� �d�Ŧ
��q�}Z�� �������b�r8�ޠ������^j���z/�|{ōO�ѫ��n2���"�,��_��f��5�)�˭��r�{P ��U��֯�I���,R����u�L[7����L�n:�����2�rD^#oe��[�b�_���Bp_�Y� ��-1�܋�IT��f��g? ��^Mm8�3Ѣq~�z�	�ȉ��L�kM"�|�pǈ�̘�c�u���lsO�k��<(�]tw����7�#�䨀FA@,�7S{q{�l�3Fݣɢ�� ��2[����a}�4�k�:� ����6���� w�n1��lgEr^�N0�$�E� ��(�!�t6 i�tj�&no��￿0���3�h��kд)���џ�"��SZ�v���QpΈ�e��+��[�-Y ��gT wv��{z%�b�RЖ0��?�3ρ��q�)���IXgh?�-�������Ί�c@�J���0�9RLG�60Bh�@�N�:!?�Fq@ E���l�j�F�&����mO�Q��n��XP%��2��4�����Vf;I��f���zS��>��*��k���tT$�ְI&#g�1w�a�^]X�hrI�E��l?�` ��;F���+��ߊ��Ǐ�o�����w�����E��P>��^Rg6P���_�����R<U��ll���y|Mo"�n�t�ŋx{�B!M�eo�[�_O��D	#E�����郬��;#�鶞=Я�+��ڕ��~��+�܆ԱGR:��;��#�;*2a���2�V)z�#TjT�P?����9(Gv�e(m ��h�٨�e6U~�Ҥ�@Xn�*��u�9S:D�-��B �@P�,l�Me�[�bm��#-{[r$%#�Cx<�]\\WE3�<���ϱ&^��k��Ӝ���=ï1�k	�k?�~�P�1[�N����������3����8�*��W�ԫ�I��/��:z�8,P�{�[x*�x��9���������@珸�w=�͎��!�4��K�@���`�V�mx�s=�,�u��jt`^����H��y϶�
[��1�J���o�� �:ׄ Ir����K�����cj?�[e{��m<�pj32�^u��|ҩ	����.���5��.t��;ޏ�a k
,�o E}���AԊE���*��{�d�~y��/^�K��1�M�ܲ)����=�,�@�l��7ht�a�}.�s���Bq�%N�)`���ȷq��B��Qd�Ӥ�*ӿ�Fqơ�3s��H:�(��L��H,g �
�j<q����9p��̌����e��L 9'@��[.�_f���X�����y�M!QE/��${��q9�+k2�_��M���v? [�� �|�1M��R����G��ͱ�[�Q��)0���lr��3!�!f^�
U�Y��H��E�m�e��ƖN��Y�|]4�@ e���f.�̒H��WZ��:@�*�c"�Q+Lj�O̡�����\���W�;���u��Id|z�Sx��c�Q$Ю^n����|�i��c�9��d# �⊰h�R8�������̕�	ӕ.�bb+�=�V��э<y���M4�l�y8��24����E����b�*[DQ�ڍGP���,��OP��P�FVU1����"����J���s(��}�NV��X�#O���}0v�5��QaK�n�`�)�C)h2o��GgPJ���B�h��O���%�$8t!�$8����R�@��!Z��,��EL7�*W.Ǖ� ��C�� ,IL5-&��'$@��VT�҈���/v���(�0�r �z��v��4)�o�:1M��l��?���L������5�s�=��Rs
�\$�N%�S6�Wj[�+�(1�Sv\3��Cɾ�w=K�꘡�l�7�x�)�D��*BQ�挵u����z��G����ou$�QWk��P̬�z��̞�A�����|5|�/lŭ�M�����!:��'��[p�7�sg����Δ�w� IN2S~�ĳ�-����;RR�gvU�\$vQ����q���u����|!�94NT�~�ήk1+;���qCm�:���u���ޣ?m&��F|�zpY�}=���'��3�i��"%�wdhi	@��rWttQrUQh}��N)||F���Q@��j���kV@D��,�&�Tp�u�"�6r����� �rKuT A�*�eCZAn@!wZ�������5��ґ~v.̄1�<�yc���Ռ����f�� �8t��5D�
x�2�p>f@ I�O���4���a��������P�G���Y
������nHȁ���� �Z�Go�Ǐ�>7`���������Ǥ���R�ed��a�=��y�]�[� $1���	��$�y�?=���|�6���G��_�� 
FJ��R��KE�����w
lT5핆�= ��?����F�zr�����u���O�l@��e��U럴�G����hHK��R���� ��Ӎӡ�Σ���#����� ��*���2��?]Ǐ�q6������R���*	�7�׽����gFX0t%DB����0��� ��v���c�N�y��-��#QѤ^]���QS	�p߮�7@����B�l��!�h���	Y|����{���E}�J=:�%��=� I��{��$z��^��Q����`��f0�=��}���뜳�Yk�_�g��A`��ӁK\��w��YeI��3�$~�?h�=x��ω��0������;��~{��mr���?�Ib�L�߲����m�[-�C	Ђ�	$~�%����N����#ߣF�}}��{�E�)��"L�U;����|���?���З��֗�9�����S(����6+�z�p��2D�k���-brD�'t��^=��zDC�aq�3l�WVO�@;s����0N�~��*9��|�A��8�·�~�)P��������	��uV��Hl_+�$�������|��=�8~܉���������N|�o?��ʷ�>�H�;�|�0�f�B+�a�wb>=S���Be��c3&������l�G��r��̏Y�����WG�9�_[7Ǥ�< �$އ�������ړ��D^z]����̰�3%U�..8�/_�k�y����t8r& ��� �\�3vr�w�՝nd����[��L�]r��OM�2�@߬��?����!��y��\c�"�:��.z��S������^�\�
wS�s��4#�� �ς�Kp>�Nv
���PS%�?���,�<�ͼ�*(C�*+FW�hy���X5�6,4͒xJ�%|�xa(J�>�
�.�s3���!ϖ��_*���u"���@�~��:J�J��M�ӑÅ����Lbw�5Q 6��X\z�;�8/�+�ޤ�������:ݩ8�?��%�����2~����:�3��l_-��G��_���7�����G����(gKKg��WX�����J< �t/���G �ޢ�T��AÚϞ���}�汆�K���=�)L�Z���V���\
���� �}���q�aF4��%�>�����Wnϧ�6�P�3Ee��~�jAȸ뇺�!p�6x9���t����)/O���d�8�����4��j0t��VYPq�a�>���a�0)�U!+�����**�E�$\|8��X�U�����'И�O��|,����yE�4����`� =��.���Qotxҧ���o(���ǯd<-��r��Zn�I;Hӥ��ಚ�;�e�\���!�"{���P�0U��|>����r���;��~��E�O�U!��X��Q�A
�s]��R�+����L���R���]��z��	�Av��Cy��>���&�[#���p��p(�WD/OQ�~��쒐���ɭZ?�vOGE���'G�Wh[v�mk,8g���6�_�BLSO7�ޒ��1���k
>�nP�_u�(ly����8�7vG6��l̈́�����K5xi��gU�3���ߺSN9���0��%kdL�J������[�|���%�֣��)�(��v����P'K�N]�����c@1v���肠g�����1H��>2��'��|J�R���zO�z�w���и�[7��m*��q�����ԍO��BE�-`�.�1�u��=�T���^)��n��Ñ0-����ۍ��B�����f[5w�Q���`˅�{�r��$�T�,���9 (Ye�V�A����Z�n/Х�11J]�]���ol��(̗鬖���0�sdX��]�J(��\~'�8�I�{��qݻ�k�P��s44�S���'�ouL!c��"�n��}V��[�
��2���,�T��>~�Ej���\��D����w�LeN�鑑K#_
��c�$�X�	K�!�̱44�f�_����}�����Ǘٹ�L��[�#�f�&< G������	�� hA���kT�3cc:�X�`e7I���=����M>�E��lZ���ȏ�TF�]��ϼ���?Uu��GEX,2��#��?a��v��c�~D���{TI�ø��r�hq@7ɀ���/����Np�O������)5[U��E�ű�j2�(��ӆ���;�ʦw��P$2	#~�En�D1�L�n�)��|ن�2�o�|��@g3�F!�\���@%Z��!�;�*Gr%+/0�$�g�ϐˈ��۵֡�7����rd�0�+W���=�[�n���X,r�|	������XC�Y���ȣG	��	��ܥ�Ȟ/��r�&pqv���[n+��ͷ�������B����e}q�.S�B� �hE��|�$;9qG�6�&��Q�e�5#9��F�G2w{�Wc�H�Z'�����L��F1�ʦ�p�u%K��-�@������:l��;Ё�h��:��d���z���h�^e>蘽�<uS�k��-.^<������Q��q��YG_$���x&�ͽ��R|�W!��6!远����ڄ�x��J��~�������De^��4/�m�Cp�MF��.��'F|�xP;�:/�;9���qWmWIU҉uF��z��k{�kv�$1���mA qӤ~���e3rd#9��f����V��|=�����O�~���e돡�{�r�N�����l�D5�T����"#�٬��dv���^y�\ � ���ܿQj�b�:Se0���N|�%����l�� �)X����Led��zNC]/��>�����~u���^���N��jt��d��Ѕz3���+t$w�ɞ�	�t�?�I�ߤ�-�Tpb�,� .�c��7c��!C�iH0 �"�b�2��t�����Y��I�d�_�Ž���=��Z�q�ç�Dl]�L����w�I����K�
����Aٍ{N3'��i����!���/�>���&BmC�\�zS��e�U��/��aD���N�4�$�f����?�!uU�T�~%{pT
�fѲ�H|C*sh�<���vo����H	��y��_�#,��"��y�������X�kҥ�_��픯4Uc/b�v��9�y�"4�Oo��%�6�$���Y��6f��l�菿,�~Ş�.��"-���!���d�_�`4�K�"��٬E��`�)d�~��o�)>�ޡ�6��<�N�؁�����7��*:ɕ�ZEי������t��OO{�f�dy��fcl����
�]�����9ɕ�U?Y��J��a��jGG�b�ђ,+�	����9��%Ó/Q�nC����=�"Ȍ�_�=�5>��%�?R� ���洫���V�Tf��������k���s���A����+�5bf�-ٯ
��e�R���8��J�|ȕ����PĒ�;��ek�q��x���ջ��4+]wj���q�����X�]=��ޗ�{?�,�������*#)i��n}�q�G��#�&uE [=���m���ג�>'�J�V�F�Y��o���̌8�,o�8�{t��ipȓ 4�S�_?$fo���m����U��M��`e�x^X�h��t��{�~��~TT��ҫM��wsZf�8Td׀�-XZv�t�����ˮpp?7�da
�>���b�}�J�x���qItv�r��S�L+ͣ�6�,Q��I�0߱0P���G������588w���v��}���\���_��I�g/d����g�$���	�j���}����</�KHv1��u�u3*t~4�(xy���M���2?qs9����ɩqN	��7 4�4)B;3��j?�86l/�8�z�!�X����SM�לF��K]ٌ��l<�E5�*�����݋,I����m\������u��H(�C}���8(��e;�ȑ��$<�&T�6J:A�OyM[��h�[Z����H�H1��#]��B�+Pk�
�I)���+�0�؏����c���;=j_1�"�4Q�v�W�2`B"7$ֿ53i�<�O��o�1�و��CS �홺2�z�K_�Q� tU�Zw�X�>���/_�n��t��jt��X>N�țk���rJ����e�6�wfB���d�����b��]���]O6�;���Q�܏U�__7�J� Z�*ó7սH�;6���	�����x�Yb8�&4UIj�տ
�2s��8j?���di�5��g���������������)䞪�¥of�mK5f��*v��]/�}��`� �d�N\�Xg�P�1ZHx���k���VW�Z���`<��9�iҐm��V����B�'�k�m�+(��*,U��g�ѱ(]�a��1y���g��`����&��Ie�lJ+\b��d���܊��?��=�0�wB����G&�]?���C'�ם!ߛ�e�<I�--0����O�����wG��>�j���n���%�^�M��,�͗vqg����^��R����f��;*\F�;5�s1�2�l�}D=�ہ��~%A��6Vi�3�7�K��re���,�d~2��DW?�b��F@3�v��DiT|�7%ڛ�w@�(�_�\���Wi�Z�gm����q"LA��B�. ��7d|B�����1���@j=#P׿m��)��ve�U�b)�S�Ud\�Ĩ���DHR�s���w�.�Pg{����^������BC/�3��?U��Hg�u���o�V����n�t\!�m�m酣Xe�FU��6ѥ/���Oy�t@vvϮ/������Q�3Q�`*����gףaק�:�v���J�qU�5"�a�vA�8��=dg/����!k�2��T׋rI;xd�U�����"��Ή��"h\���uH�{�֥�Z+�0k�3]�	���� ��;e�ޟ.�X�"�џT�Q����n��B�Q��M�5q�}���L�SgqXЏ�ଡ଼�؀��~ȹ���t��&[�<aKK�if�O��Aš��,��3�o!Zu7[9��E��_{N��!�}L�{�g��q�P�]ҧ:� �(�߬�o���F���i���6�%\��,d�O�g�@�����
s�k*X�g��6����1V�1덺�J�	�?ț��;*��������؃tYDK��璁���{ZYiu#/�BOw�-�&��x��.��i���UU ݂�ۺD���La�p�j��G���y��������%�--r�OuAG�0ض���;����_��{)e���e��y����b�����bQN�3��u�>XH������䈗p�6�?�����ف�$?�@�G��he�
�%���G)��'k�`�T�{���,�Q?�`��o���ϥ��A�Pp�*y=�s�����?4D&��!�r�م�8@ƈd��5�倜yi�o ���� z��ZK�y������SC#k6�	ԅa7�zJ�r���h?�f"�9�ju=q}���$v؄�9>�0k��ٚ�!G������C��Z���iv�ߔ�kt��]g��T�S�6_1���%��
}F���dG̯�7�<�:�'���<�ud�e���.����Ժ}��rQ� c��C)�W�쳛���>}-([�#�-F]�u�����~�����<�H�_��\x9��B0g�şe^$F)����k�w/@��⩞g���R��?3�����꤁�o����NL���MY�����m3���ݟrm�����F�W�oFN�OH{�>���v>�ct��������8_%�l
�|�{^e:�f��6�ͺ(�~%���Lmߟ����=%zX�Y��H����з��U�2�.�.�[��Ew3��(S���?�t�i��A]##F_>;G�����Iu���^��g_����]?�29�p���2��IS2%?�r����@Z�*Ye�׬��!�ߜi*;���:�z5�����)���o��\�.>�zv��>L'��Ιq<�G�:�7j�+��>T1۟���&e)��C�^U˟����g3�Sa, �mtt0ՍQB<���=�w���$��>��g�Ή�{���é�#���!��V�A��d��'����^�nkʫ�<b�I���6��eRN_�7�l���C^H@��os��� "ohl���)fJW��l�_s���r9���.^[�h��,l����#��o&�`����
V��q�Y��wX���^��YEԧ���H?�=����K��xc*B<I�Ηp�R'�� 9��e~Q��2�������D�R�_/\��2����U��l����'���i�[T�^,�m2�u�=A��[�?lL�e.c)��v��f��%�C��y�"���,�M5��Ip@�� *��u���職�O�y[6	$6#�H�����H��9���_������6�x
��4��q_�'��0%nb	���6}:'}�s6�D�&����m�U�U-����2�HK����\����%�|#�$M{��G�Ԋ;tlq�\��o~����>S���\�nZɶ]l�R�k�/�b��8����y�ϥ�eFo��𖿍�&,�@>i�.[�߿��u��I����
q��O���#=���	RkPOcԈ�f=$4t.#����{�A7M�pXJ�/��OB/ʂw�m��j��e��Ză�>�)���?���*���A�<2��~Rsi0���������}�=��6��j��mqC�G2����u��@c�H���R8��&e�J�T���ϔ�-0����%o�/��T��.|Mhcp�t��1ju�_�N�8�Wa�^#l�%%*�t^Q_�����]�D*A�������s-֑�W3"���L݋�=پ��,��з�k{K.
PA�� �`ѫuv�a��ծ���Bb��è�Y��kJM1���0�͍9K� ������S��d��o�4�&���n��Rd�:N���IJ���_�9�&��k%�����/�%F%'�!Sii��3#v~�[;r��*mO^�p-�v�zf �yu�J���	���*�U�I�`�VH�_Hf�c9A��U����:��<HzӲ�P��˕PW;� �4��T6�	r�?�KBzPMd�3�$�K��w�lg�#�	[r��{w�N��<�	|�V_�
�U`�&0KQ ����ߎU ����u�֥�w��͜Ň�O��!��|I׭��R �}�)6/.n�*���$���&>����2�_Iz�|�����vc���K������l��%|5z8�]�z�_��X���*�
`��po�7���,���2H��S��+����33_�7QO��k����O"d�����z��k�Y�jeћ��53ʱ���X����κ2��%�T&�=,�ڤ����zy �R�1͒�hW��s�4m?�2�A���7s�7��Ĵ�L!%���}� �L��2d�� �ktp��r���Z����%�N��n7��7�RQ����w'���"����Nw����!s��LEA�!��N|�|ח<��i͞�)�o�[��W�OU�׸g���6�`�?��x,��#�5�Q_ݧ�v�K������l�rzL_�	@�°��Oj��|��{���?� J%z�/>I E=�ҭ	�����3C�C0}>;6�`�KY�$�[���k73��98������|98�Iψ���>����,�}�( �� ��p���7aN7Z(T��HT���(����~".�mN����A4�{t����ކΖw4��\��(
�D��F9D��	!������ܳ��h�"����fsn@�Z����(uN�hr|�QtNL�y���|�P��˸yS�N������8�^��@f&�\J��l`��[�@@�p�Z}vf����X��y��l�1��7����M�;��?W�pNwU�F��л?�3��s
�O���/q�t�>ye��遫�p�&�T ikns�V��A�c
_����x��+�z�-"�� �n���l��D�<<��O�>�L��;����*���1��ߵ�����:����s�e�ž�l�Ys�ᬬ܃���EC����t�t.��{��ڜ	�8�zH���vwٵ�!�f�F�t�.��B3��Q%�,�;�(PB"��˶����8�A]t���{ �ǏEXG�N����+}�-��L��Y���8ށ۹�nx�t4?ё��r�H�p�CF�b��33l\A��,��^��]����yw��͜�zF��&k�K�L������]c��d�V��7�0��{]b:�]mni�^�6o<���0.yU���,���r�z����
�E��ߗ����;yn�`�}���W˰���\7Ƶ=�E��X���k��`�D��1f3�2�o��u�z4�ߒI��]�2e7�Ts�J����#s���u	�~꺇�M��5�v��<R:�滞�e�X��%0i3$�Yuww���fƃ��m�yyxx�i'���{�$�W�6|�eN���|�Ž�����O���ܤmb�b�{�G������xq�g�f�Bxʗ��,�f����}�P��Un��ĥM�rwuqk9��UHAĲ�TGQt��󧼋SŔ&���S$�����<��J�xA�=�w�-�zz�1�X���"�LH'v���&Z4��\�}u˧=�:"�o�
]IT����Kd��������_d�6�Y��^����j����Z�1;�6U���P6�%O�Gm�)8>S���*��tL�r+���Hſ+Md� ��t��V+&�O�x�������B��5/�����=�cb�bF����:@��mmv�ܠF{��R�\f���l������<�XFy�$e�ZK���u����tdg���O��h�������Ugҕҵs�Q��"����Y	��k���Ňɷ��\V)���khGX�cC���{�㓁�+.Qś�}l�쓵��$+�T<�Sk�^���\Fmf,�Ǻ���B��r#�)�y�R�?������]5���%�5��xC~ʽ� �
�Y��3�O�̇+�(b)��:iLE>)�H�uom�֒�S�� �� �|S�]��왌���lQd�ׁ�&cużEII���_�,��<�֗�[�����Bt���m��6��)�GAȎ_�N�9�鉂7b�?�܍��ޣ�� x��-��Xv�t4wDT��i�Ӑ��
g���>N�ً��[Kg���fx�^�S�����%�}v_j��}0e�H��m���!��e�`������(��g�C�e:*�Ѐ�(Ώ��-��%ܟ˘�,}�?��[e8ھ;~y:\�������49��j�Mc��9JY4~�<r�Ό�L��1�Mxd$o3z�>,d�èc�Bz�`�;Oׁ99��/'���;��_����S%��R�����Xm�aHb4?(��Ծ�ƭؚH^���*JF+P�k�w�v��E��̈́p�(1� �{Dt%�����x�4�e�?UP���I�݋O��հg�P�+�M����������x�5h���ٍ�&f+�ä�S���!6�X�z�S^�Ӄ��@.�'(�����q��г�b-\���Byr�,�f�}�9�>L���zYT��H�KQfU�z`t�R�É�ٺ��cI'�h���$kP{�����J97N卓iA�0�����#�҈����߮��]����4~�h�ݕKCK�����_$���p!l���_N�ݩ��ㅡ�����n6E��!C��-=��n�6J��u�X�A�G]�7��J[5)��o�f�&I�7��G���D��r��{�R$�z�X���8�~��۪�����՟�W����Qf��)hO9��Yp�2��]Y��]X�=G��N��0�x�9��#�3Qi�XK�?�VΖ%��.U�����r&��Ǽ����W�B�c��0�[] ��'��?�����;��;l%���zup��ߖ7�䀡�j��$����xr���)�pnO��,�^�d��rW��1��b�k�<�d�p}�7[�D�l��y&u���	��b�5R�f*�+?H�c �����Y�U�FQǰ����n���y��_�0Va
�Cՙ�ŞG�`�˯C2rjm�{	�3�TI�l熷kr;N�W��r\��׸mf@d���16�# ����2��l��D��W��V�ߧ���DEI�h���8��O�z�`8.u?�j�e�j���l����f��MNKp����J�U�8CW5n����H��}۷��L�%Y��=�����^�A����sd�~��8!Z��K5&^�`�MuT�3�5����&@��B/�^I�qI쮲q��qk1{�Q�۳�+=>?*����IR���ș���Ɖ�v�W��Qi߳��@#�,�xx��-��tw�ԡ#^X���A��7ԋg���92�}��pT��[�T�0>�rT:U�D��:�@�x���������dvX��r��,�8�u�Y>�L��)lc�f��1�(��ͱ�}8	wn��Ix����Ba����T����^G�*T���"��V6�JL�,B��L&~�����u��}���((�uB������M&��tY���@5��i-��5G*׉�-ŗZ�g��y��4�	X��_.�N�����I�,���3/qG���9`���-�����A�P�u�V�S�
�3{Ą�SQ�j��z��u���b?��E��(?oBc��̵@x�{*��>�޸´�S9sT���Zq+���2�������wxr�b��n�ׇ]�T�#�j��\���X�	��|���1s�����p��O�Kú�9tA�{/�ja�5��>��q��E1H�E�W?�B��j���~>�9�U���1����	�0,�a�iZ�90i��G��H�XF���MF��e�J��
{�z,}��+]GdH-���᧳9DD�11WUL1�^T�p��T�	��(�s��>t`�_w/9fI���PT[TF�Y�7'��y�G�~e��� �M'|��n��-�po�O¦�����@�"is�B��;��O|�W��%�JKߣ-���u���F�F)��jg���s����2�S�s	h�x\u��닻�d�9�2����.1��O�++n�s��#n&9��0���F9:�t�6�/����0S;^��/��}A"P� �ih�:�5K��&W�4�/�r_�t����`ޱ�Ha�1�O"�~'�*D�,L9�9�0�{����߃�m�N�H����4��yZ��k7�n!��-�mR�u\�i�Q��'Y���잒u H:�Lsm@&�[4��I��CS[3HK�W�2��s�I�6m���L�\&�9x�+imGn:������G����w��(7G����������d .��ʨ�I�˳'����C%�[)0�W�tD�|��3+��dU�!�R�X͗C��#9ÓBj����ߙ��^��X\�T���^ZBb@���^�8��ޤ}&�����EN�,�9H&K2��K��~��|j�Wϐ5�7Yf9h�vt9x�EU}����4�đs�6��C�>��h��{ک�p��x\b���_(u�r���Ds��i��؋Dg���)ڡQ�v]Ij��U-���|G��uc�n��挸��h��ٛD��y�K�i�>}9W����r�ں���zC��-�J�FQ�������+��o_dg�p�v~�7K`�47{5�����`��WhD��0�4��Ѡ����;G
��)��«98�~2�
���V�_���`��X�����"��+��[&}��_bb��X�3�m����a�+����:��&j��'M�n��;J)�����d�~!���G��i��b�7�#0$� ��N��NX�E>�/�k�c���:Դ���S|m���2�؅�߈ʉQ����%�7/��F��{?��?��9�)CT΋@d�8O�����L妊K"��Z�B�+#'BID�G&X��i��{�T�����ȇ��ϓ9�4P�H��ί���*�p<l�g�T����)(���K>�q��0d������a� ��-���x��i�V���^��GDЫg�T�ؼ�i@MdeE�����;Ŕi�K�a�+�B�+<J9�ᬬ�	י�&��-����U�J�����9�)�]�L�������4�b�Kצ�e�b"�fs!l�D�,e����n��T0ƛ��:wA髨\M���~���J���9z���w���%��|�~yH���������wK�ے#X���W�6'�I��H���fց��~r�S����LԾv�43/4⡲��2�(��D�Wa����Wp(�����=��h�H�ؤALP��T� 3�#d�c�+u댾:<�Y���5؃��c�ǔ�0/�Z�fP�kN4z�e��)�6@ؤq��j� ����-'��x8\�ߢ��f{�J7�Wa:**�q5Ùq��j4F�O).�ĕفI0��<��u��!t�y�7��ג��x�l���*.��![ya�?n������2;��)qZ�W�~owV��2S*z�a�AD�W�Q�9��ؘ1[�]��[_m��\Z�rܡASb<I���P��@�M�@ćfy��jJ�gf��N�+_o.�I�	i�'�P\q�ƸE|$�+�i�� ā�����:��B��t~�����qa�)���)����,q���'�0ע>!� O�8!������T��ǁJ��R�2TIT���pu��Y�~�h�
zh��Kz�`�辖��J6�Q���,`��X�zn~S��w�*��$)^,Wu��߷%����T�'b�+:�����v��r�蜈�yW���������X�Q��\lL!	i����+��FL�3�l2�A@:� �s��o��9�����DHα'��I����V���(��������E�^���[1�C��·��U&t���D�6��'�jL���;��{ {2,��>'��#L���M�B��@I8o��,��1 ���>����<ܗP�qɖv�����*81i)�$;k%y+1𫿥�.��K�����\�g�� ����B%e#Ϊ1�sβ}{?�z`�b�R����xu��_h����5N�X<&=���1���\�tq�w�G���{g�f�׬x�$$��%t9����wuz��F)b�~���H�%��)ds���?�+�]\�. t�'�x7�d�8�?]7�!C�դֆ`o��T���4�n3�>�F�����z%8--�[��Q�YCa~$R����HY��p�p�۩\�t�w)�?�;��e��ϖ�)`���a8��Z [��@��Ṇh ݱv��JJn�F��_��:o��稂,�J,X9p���6�1KK���鍺z_���������Z�Ą���u+�:Ja��TN��d������!��������V��:��w�0Q<˓K�	n�x���21������\�A�2P%=�'�l̷��I*�D%l�����Y�)���_�A���%��4�%�d�B�3�&��9F�D�T~�[��)P�.>�j�Q=���S<��Z�(ޮS"'��ď��Aa E��-�k�	�9��E�/JB&|�_5�TG�Z���?!u���	^t��Z�y�xF�y	O�x�)h�������ɤ�M�P7Qo�
a2�H������.�<%��C��X~��S:�����p�7�i�y!�n���kb�u���i��,�3Jܵ[R��]��D���k
w���y�;-�H��h�;=��P���˒RY�D�q�vّ��w�פPEL�Kz��$է^��d�͈���|�s�jf=?����9M���ů�W[m�3���͛0�7�	:Moߒ��7Ͳ��3c���}�&�xmͨ�HS�'<�ܭF��!w�	ӵ�zw��̚�g�aafO��(���(����|Z* �^31�vsv�S����
0#��A݉��;��MW�������N$�f��HT i8��6��=Mzs������o?XS�u������=���XC��~q%�$7�	2���s^]�<�N��XN�4�� m���1��l�p�p�&������7U0M%sBݯ��U~�IK��O��#Z�SXҢI�%*�(�e�/��F��߅b�fm0颀���+^��;_�+^��+m����B�x�-�>8;r\�f7%=#���j�1r��ԒeJzp�m�:�L��!�_�0��������T�gѣ_e�������s�����yWHmȆ:����|y�M���V.���H��PG�فN����$0�?+ f|�Aݹ�c�N.�~7���#����J��r����8T��(�\]�$ �t�Gμ"T*0c�!NG�a_(����J��3w����T
���� U� �[$&�AE�G�Є��+����?������HX��A"|���73j��`^js_̏B�s�����S�.
�������'�� ��x��<=@��%�e��ⵝ�M�9�iczB8�l�
b݆1���y҈J͒��tA�ܻ�,/���q�C���w��͈�H��g��Gv���T���HH�1s03]�23�#�Ev��;/^^Yx�-�Q��[�f�5�x���ò���w��Z�y���L���O]�:��>k�6���3���n�ڱ
'��qt���<y'<Mz^s֛vm�6��nr��M̙�W��*[|*('��d��x�Χ'R�$?���k�SA�&7p@��Y����bà�U`���y�U�Q� �!M}����\��5Kc	����$���|��wDu����3`8�ՠ���D�"|�����
�>��^�����Җc�! pxl�
��s���	�-�G�����tY+�i]Y��m/� ����P���\�5`�7�RL}���� ��2�i�f*D�a�
�̒�:7GrD|����O���e�δ�@8�\-��i��l��i#�I��M�p�,ñ"f(RQ�Ж<�$�cP{�	���'����3��N�b6`� &��Ӣ\;Z����&���������e~�x=����>=¦���PG�؛@9/C�y�?�zu�9�I'_d.�==�i�T�����'7�ٱ�9gat7Q�F�/��	������IqK�E�>6q��[M1Mv'��P�*����\���}5���H���mg��k�0'�47�m�ycF��ಠ��N� �?�b}s��!/��{�q|��-o�)�Y���:��Fr�m���F��֐�J�����y:^�Lw[ăO�����3��rv��~+ Lͭ�����y;ZI��~�����Z������ȹt�08�ϫ�c���&�tY��Yw2W-bUB�5:�C��'|�����F���7z�
��In�|ߵp��<W��,~��������_���I�F���\�ID�"R 	4�H0����o��zu��s�!FF�	iD6�j��i(c������<+��+_�s�*�����Ȍ�YhKp��ZH���RHmG3�P�ؐۡf4xTa�=�D���F�]\}���n�1�^k��Q%�=�ᑡ�S(��X��-������X�Rf�e\��D4�����]���I�
_�B��n�8�N_O��W�fgI^�`A�~�d����h��w��Z�|=�y�&6ݺ��^�����Լ��W۴�;
׹�w�]r�U?�����]~�� @⭿;Q�,|�f�:Z����� K�s�>9ϐ���~Gf�
�	C��}R�.х�Fq>l��z~g�3?$;`���1���F���;f)U���[��%,2d����g��t�����O1��5�����m�)q��hw4��X0�F�	�����5{��`�!C�~�;2rOR%���)��C��zB��}�di���Ϡ��/�eg�����<X����	;kତ��s>rI��n��2H�����mf��3�\�r��P��d������/��|�Ƈ2�Q���[9��@<�s�mw�_�os����+y�7�ϓ��j���q�����)�[�#��A���@u�bOy>�,�X�IC�޻�w�7���KY���W��z��o�2!]�E=._mG��䌰=RzAh�u��&���$����t8��W����w	d�����<͊"��v��f�����\���pq�h��Ne�I�<�b.����҂�נ���3�Ƨ��C/!����bD�#����O҄�%�/\e3����[�?�"�n��ϕj�)������	Kh3��w���h��=��������핖=,�{����h��"P�ܭ�%�u�����n��H?���
<�M�<5�z]f58��/}��|�2�6K�a/O�ڤ�������| r��Ǧ.�e\ӵċ��!�3������6��ؚ"i����n3�s�ɷ���vX� F�O���V��N�l����r����W�x����2�:�z�a/�Z�G���S54��}-�-��L��^���_�S<2=�A���+�r>���n��w)!���ṭ��ԙ5�̨��^��b"ꗐ�6�j��MA���=7l�M�s�g��-��n�gޖn����0��w��Fʣ���!Z���&׭���З�}����+�WDY�7�t�&��Ǘa��������g�+O�p�/���/]DZ��#sl�����俊���}��E�X��K?�����橚봋��K�ŶߔyZn��LZ���B4��g(����I?��r4��V�@���������C��h}�0��{�����W"v����<J�Z3�rKv��9i�c��Bg�9b[��٦�f��H&�V�������?^"�@ ��	2ұfy*Ը�Z��j�E"� �O�+t��J	(��6�E0џ�jY��s�S��A�~k�3^i�
���!���,`�}>윘��2*�1��l�O"K�|�;u�������Ս����}�W�(�'��r��&tZ
��*Cճڸ���Xo|6��sq��i\�v.�VI,�`y�o����zn�ş���� �g.���g++қ��ף���a�����˟�yB�.}n?�cv׊�m٪��+��-	�N��$ 	����< Ҍ��8%Eh������O_����*��` *��HK�(�ni����k --�C�Jo�6�F�9�g�����^O�s����tAmzM`�.����߫*�`�<y���+;�aj��Q��ٶ���v
�_.�l�����Q��o�af!�����PpǏgN��Bg+�c@�T���*�[��dD�A���7�_E����.*p_���E���ˉ~'�t:ț��nޱ<��[NK��C4E�n�x��(��FHլ�k�+F�iF�U��\$f/�^����������|]~KDD��X�"��ۧ���,UEYY���x gԲ��u��&K������#qu�V��:x'F�Zm�Z�����"�j͠��	��zy>a�r��,����dq��@�� ��gڅz�N��Vl
\���$i��@���0Y�º �c#>�~�4�x�!�ْ�?�y"wI(����!ZI����t� 655:G����Ҫ(������������1��z�����O�m֝�0��.9w�+b��˫'��~3My
|��0��"���N:Y���=&o�z�����V����
/Mj���ߛxb3(^	"�VM� �}��֐�c���e���o�[jF���f~3E��˙���`0z��y@�b:H%s�W�DФ{߮�������EK{�4����d�v���#?o�3�%��fWNn٨`���a(2�b�:� ��/��C��n�'��I���7?겯$'���DE/�S� a!b#u��fH�L�.����+�R_FT��b]��]bb�����kǯ�.y�IZ(��.94��Wn�x�m���QM�AX8������u�
��O�]����8}�blNF��1�����Ǿ(E1���_�T�3�
��-�t��+[�}�x9�nk�>����*萇~8]�Bв� ³��ڡS��z��PCCK�C@��G���ad�V[��dF�b��h�`i�C�+Yo�*�qsa�������o���3�A$����]�+����3��7���������S/�.	�VgKw�{��j*J�^l�*��N�u��bl�K�PΎyV�������EG���&k�s����=�p�\d[�8�H2�#'�m�s����ٌتkJ�z��R�<�?�~[��u����V�G���9��o] ��򖓿`d퀂!޾"8Fܥ����G�$PP�4-?Z)��o �[�I�T��(��1P����FEn:ı�
z�̟����#��	ߕ�N�V0U+bg���[���#���~K���3�|pE���R74�-̿���o�
���'@;yX[�t/���'�ܒ��Zl(9��Xb!��е���(�*^ǑYb:2��Q�~t���9p�B�~�o����O��\��x��>�Ou7�_��onwP������Ќ�޵�0?��JͭƱ��T�WF
��G-c�o����@D/���:�Շx��@���%�l��:��i������a}�g����iwΈ����L���z���Tg���a�ϸ����?ToL�6'h�6_�|����\�C�7�h�7S��V�p:���/�p��jH�.-#;(�R/��^*���f��h5'��M�ǻ�i����\#6c�(%��ůGKȤXx� 	C
Y?��dп�C�t���鑛/ħ��Z1Ű��m�.�nXB�fqbM[�����_�#��&�i�g��V�J?.}#3 /"��J����CJ�熺����E�㟙���-2�����'�(��:Q?,%�@K�#���]˶p֎O7��H���'w����2K�ӽ|�_��#�_��ϥz�V2��OIF��T��:�})	���⚡��E;�5k%`wu��`x��6�y������r}mAozQ�p���F���k�ҭ�L����V3!HZn�����'.Hۈ���T��`��3��3�%u���^ﵷ�"V���t\�����]͍ۤ�jZ@7~���FP��$
�Y���� �6I�j��8O�3�E��pわC;��H��N��# B��x?8ϸZh$u[��n0��u��P�j7�����g~u{
T�VU�!��ŉ��X���{R�:X�W$�vn������jT�I)�c��R� ��K�j���X\j�:���ĩ�NXN���h=�rr?�!��:��QJbO.K��gZW��U�.�b��i殓r���aǞ^V���}jn�w�e�Z���5��bN�B�lGf�Dȁ2<ULDAp��ʒ��2�_��d�8���>��~�H�l���9�����|��}�Te�<� ט��I�JJsj�%s�Ԯ�/T�:2�ɞKV�l������q��N�/�4̼;�����;'��:�3Ά|��X����*L��ba�[��޿�O��3�a����D7��^� �����s`G��&߿o+��hv�r&�&�WhPn�	���v^q�ʾ�u??f��G$5��014�t:d���M�)n��Zаd�iay��bO��E�6�ƴ0�v(��o�����QSOG��=#�jĠM�֑��\���=���#�Ux��e��l���s=��I��&|��ߩ��W&�\�w2�nC�������u� ����ӑ��|wi%�-O��ÒMO���SG�E��p�	VlE��jv�Mi����5�;sIr
����5�)�f�j�����_�GK�f]��PǿMn9r=���t�����tW�JK���-{��:�D{bV�ڂ�n�������})k�{\�i�:? ?�2�#|_�/�'"��Σ��3=w�S^H�J���E`]O<z��V�x���k�_�?�:@Jļ��u>���+wb�S���1n��[��/mo���b�3��Y��7�pu��o��ټT�����	8�@�|j��@�<��`�k�ʉ����,+�%݃�,̜�p�O�n9�u#�����j��h��6*2MHU��� E)�T� ��mb#����h�w��=��=�4�k��o�_["���A��T9�OZ���yed����8쾚5]�7�j�bBԕ�;��Vs�֏��6ϴ��[��U����p �4��4������`�z�=<v��l>��=��7��"lccc���˗6+�����$��ɘ����;�����������M�נϸ:�}�D��VW��s���@��-1�����!��B��t�f�jW�;�y۸��28�F{���
��ѕ�S|�rrko~����jx�pD~�i�Q)eے�����̷9Ȏ8UUm�Mы_X1@��t~���=Xd8 �gd�= �Jw��=*���3�Ez�1{�jIb8�ɣ�sKI��(��j˞����\��A�lВV���5��n+����J�����n�Q	��drT�ȦK��Q�=8L�O�)����"�T(!�+"�p\5��%�����])%%�=*NM[;����p��]�����k��b�y+"#s��߸L#��Z4!��	$'��Qc���C�:ס���_o
��)�|��6�og�"�&���t]%�}.l�D>��7ū���t�-���-��A����B����z�}��Ow�WUUuj?��}���w<Oi+$���%g�2�%��,�h�\�dI��O�N��?¯����sޘK̋��G��!󍅘4zA��'�$fue�\��̳�qЅۓ%G�v`��wW�Y!8y�[��?�G \4aD~nZ�v����A������L�"_�M�C�b�Hz�c"W����_�%�z���a�R�7��-3*��WO� C9�����GU�)�C�Q�dvg#����f����ֺ~��� Lm��K�W7�5���f��|8كi:��l)GAZV�����h˷Z����M3O�s��5'y���\���|��Ӥ��ׯ\��*�������/����I� � �&2�����j�	����^�vXLFd(��ǈ��OR=���@�$1�h���R��=7.���.Ӆ�Hh,�֣��xy�Y��u���Z�9LA3�3�t��yP��q���{L�Fʹ*�E҇�o �S.������)��ӨT3�_��s�9��{���s�4+�F
� �4}�0��9�r"cN��#:M����;��(�Y�+�(X��c؆3���!�t��8���YJ:�=��C�9a�_kEA�;���{mt�O;�93�cX�k���m=�r.}Y��א\~p�x�kL�뾝d���Z���T�������vA�o�*f���v�h+�r�Q��
'������M�^Iy��c��!�I��z�N�KLni���L�_��R�"or�e�!L��&�|���Z��L`cR�Qc�7R�t<@� Evt�VW*JM$+W�LPA�S;KX4�0���<��Cs��Z�g�xnqo#�� U�ԃ������u��y�;a��M�X؄�y��KT��0��If8s��ϯA9��[g+5�{sSN�n��K��.��*���^�����(O�0��i����ym �}?]"m�ի������I!������%���+�>�C���a��orF�����Q�p�g��Y�ټ*�˙��4n�D�|
#�o�f'�ڦ �������}���}�vn>�tpY�Қ9�;��Ff�hbd�7���i<���&���3,K�<�@ȑ��i��m�E~Z��k.��js� �.�Զ�CP������9_v���9-@�5��TOǘj��o/�~I��ʕ�ʔ��U6�S4�����sw���UQ���/��:>,�����Vx�Ը�N ]�G
~2,Fu[x|��IDDΕT��^�X�+.��B�6�c���.ro<�I��l��k<6�A�oK��V�Sh�v�R?y���6�;^�xci��(�ް��� 0�ɗ�F!Gy� ����8(K�(q��o�����7j�y�iﴟ����zFᓵ▂�Դy%|�<]����i=w�2���\>�3�<�J���@��,�YN#d���=qI݋�x�Ku��|0����9��B�L^j���Rj��uU�k�p�"h����R�4x�)�*�Ͽ��vG�9�(K�U��s�͑���<��:b�� �ӌ'�Gj�=��>�~��}�����ˆۏ��?b��A���z+�πyNf/�-�W�9&�?��k����ɗ���l�Q������<�A\t�= h��9�oz����(��(R�xuY�$��H==��b�Zã���}����r66���ll���=j�ӄsH���8,�����))i`wj��J��m�����u��Ȯ{nZ�OsBio�t����6I��+�=��|R���֏�J�<��_��aW^�5�~�ֵ+X�>1G݊A֕_�2}�U�͍�H4g���:zG�Q3�ǈ�G����< ����8�}1-�\y7n�4s�G���n����Ժe" oS�	3'�*�PD�������L�$;1���!w�z�6���k1!�)���{�%`��~��r��V�ǿ��>ڣaZe��^:0�jh,�}P�ԙ)��P`�̃>͕��X����92����efQU a�@��������!!$��b���L�e�
�>͇���'/�ǸU7�FT��ݒ9��p
X�oȺ�Ԧ@r��N�K�b�����g)�pT y��Ƞ��>�́��;�"SC1�ᚣ�_ZLNL�����H�`U�ɨw��j��φqD1�1ɬ2���S�O� Z5����G�n�8�ؼ������@�J)m�[�!ڊ��[�BP�+Lɟ"Cx��@V���@*ťףZ(� �`�����;���ѓ̳p����4~\�r�|��qE�ݙ�Z3��X�����aj�aw�U�2y������u�-�u�Z>��B�1ͮ,*�}G�~���e��o����|�\!�ƕ�4v�O��ú �o��WN�Ѥ�
��"x06ڬ�f���-+�B�\7���gejM6#�d|��&���J�x�i�u.��=X�t�JB$6��v:�&����JWw0+"����)�����$��=��Uw�
��z�y3�p+A�%�d1��\Ǻ�|�mi�"9p�W�,8�+͘�-�EC���+��%xΒ�_km|�!���]����jBr�v,`a:'ǃ9�f�)��2S�5`m��9�,7m�{�[�o��{�,~OA[MG[���yC5PT�ќP��:�?���b����eFig��.��b^��HU�)�=y�餽~KB�iH�@$6_<դ��2�^��RZ�w��k�{{����ki��g���[j��z�=���D����>���i�ekH>���K:�u-K��ۆ>5^�����b�������uh_q���l�!�����B���; � ں����0θ˟%��ȈT�?���m�		|k:V݅�h��Y���*�a��9��*�&k����c�/}fĹS�<({�����q�DMo0CVKEUs_�c�tz'w:��I�E�T\&W=D- ����e1�E�f��u&��P���֍A���50;�R��?��`�}g���Sr �������?pp�����W��ٻ=����'����K�y^�	��
��K��v�ù���=�\����R�������00�0���M�������ՂO��z���ټg6�x��-�J}����2
T�N�:�P��5�sUXv���)3o�ܪ~� O��pd�B<,��͹�w���j��q���v�A��37��C�ό͗h�v���rD���
��C����X>;	����cSݢI�z�9a���%�ց�7O!<�2E���Ca�X} �}i1�l�0�{��Ǝb���x�$�!���w���k�(p$���3Ȏ�zJ%R����͜*�����0K���U�^�	�B�8�{��$��QQn�)���a�<<�<42n0,����
H�coO�� ��Z�qk�pV��%ݗܲG?pC
��T�'k�����#�N�c���@���+��%�e�S��K����{��=��m��\d�כNM�X��M�����S6���o\��'�2 tIT�}���I���ƫ�������0p�k�������"�\�sT�Ω��z&G�����a{�q_����7'%I��U_Y^_����2%9z�Kϐ����i���6���P�E\
���$c��"�Z�8%e����YN�s�ʮc�8�����?��׻���Z�D�>��xq7IH�dhQ9ݕ|'����X��]o݌IH�A�����p�������M�&%��t��e�Ic0�|�a���7g��������OMu]�}���ҿ�ٳ,Z�燵Ɂ+mv�<$$�T�eS��gZ�h">*8;d@B2O	�I�,u�����ʿQH��/�]ל�D���,7%vX���#�N�W�fsuf�{�U�;�h.��aF��C}h_TZ*�Lz���e��
�q�6"zu%�!;|�}[IK+
sU���7�z
U��­��AG�V˿����Q�P�N���iL��S�􋊄�� �60'���������Df����٤��ey�M9��@�@�I۶��hUǇ����^��g�Ƕ9�I8��E.�~�w��PX�w{3(ޔE��|l3�;������&̌�i���P��mE�m�T���t~1s�J�f�ϟO��u�Q3�*E��j7��߇�r6�=|')JGZ��?��QE'3 �0_�|��Q"���Ci3�FǙi�������qך M3���#��&�TM��@<�Wz�Q��`��00����������	II{T��	+)i��@j�́[�[��4牦f�~Xm`l��d��,�7t1xqDD�˪ܖ`-��L��������(�E�� e�ق.���D�����+�1[P���I���f�P�	��!��J:^�)jG-�&%y�dP~�[8�3���bB��Z_D�+���0鰮{�o}'����$$���h�~LD/�=M��y���v���^6���O���jTƦ���F	���K T�X����g.�M������"o]�%��
~
Qf�o���>9k�W��?��<���oV7pq_�9Gh�A�t�NN.Lr�il��Nr���B�ؙ�.�L�j���:�"*������+M����&R%�N���a�F�:�r�9�}y{��d���n���_!	�@JK�p�8�Ͱ�å� ��(;�Wx;�� ��0w-��{��@�/A��P��gM���L�����$b�^sG����t������s�@؂C��-҇~��a��|@�ၢhظ��Y/u)cb\*W0(��'�dJ��$j]�v����<�e�%��dP�ZԜ
P��A��۷^���&ZT��˗�����и�V�h&!f`VE*���*����܀���J�S�ݹN�?ΚJ���0+��a�WP�U����f�5p��V("U6�spH'Z�ќ$(J ��"�t^�NU�Db�� �E���Uzu���g�ZT��1�;?a�lD��QG�άO�`R�k��/d�J�0���ŷyyy������gZ�M�0�I��pޖ-!p�3�:pP@0��-8$����pK���;yhXs
 wc����3B����o���kc�i�{O�60��:���| z����N'Z4��ŬBg7R��V��r�HqC���unn��j��)9�ܗ35�4��=�j�y���
��鐭;7"6�`��eP��<��ymZ?r#ʇ�������kh���u�k.��c�1���V��'����rn�� y��j���A�EFą�ݾɻ�9pf��7 ݄��8��U���p��*��O_I�򒁁��^8�[� ���EؓEXI�~"Bɿ'��O\X�˦b���[J���1���b�zI�O�2)2��@d�OG���u���!{�"y���{�1��1�̂�:�7�7���A�U��I>ߧE�ܻ���%�/r���
�q��ai�A�,��{� ���B�
�}�\���ý2���$W��@�W�E>�`C�׀G�	�}���.2�S��V�O��K�;���F*^ _�Tu[����U�M� )�Ϭŷf����>�ې����;��D.r�>I�(�ؤ5W��������Z>�����p��i`���>��S5�Z�4�½)���Df��t@q�XʹU�6��z22����ػ�~DO�A@��*$�_��Ds9��M��P��-quz��j��� GmF��ʧ���M����� _U��vk�<�����s�	0ǽ!����b=B]��?>�<͆�$��Q3k��l�"`���JT�'uZ��@�&X���c�[�R��r�Jk7�@�<��"d�֚Ĺ>������1��;�_<l>r���ϋΞU�7B���7:��O!K�1���y�9�^F?�.پl��7ֽ��b�%չ�������|�I5-0i�QkI�;���{u�f���cR�юm�tk��Qz��Z=�+�*P�f��C,*�%p\��{��$7�O��R_(C4b��AUk�Q�Ps�4W4�G���^�8���Ho~U(擿PߩV�_W+��/�O�G>K+s���R���L��;��]/�j	e��OM�_N,�)J��f��
zi�F��G/�h��v�A����)���ѵ�ʭ2*�qW	f��+����tP�򿉮�5����UqZ�<���5?j&��'�WN�Hq�~U���bO�,t5gB@���������#�Ѽ���;` E���nƹ(EO��5�ѣ4L]�;����$��5ӱ'��$�h.��&f�� uT�L�����S��@M��+|�[����~�XHJ-�w��6�R�G��V�5�z|N)J�U Us���^�ε�]�3&Z[��h.rS%bw�=n�����V%���A��-�hH[-]a	6h\��^��6ݜ0%j�4��8��X�~oP�J*�QЌ�v�kf�MQB��Ƴ\}���� �Q���R&��> ��5H�gY��oY��$y��,XKô�f��-gա*c)�Mۢ'�O0��-�o�0vr�����D�ʛ�8b��um<k :�iQ�s�{Ό��R1I�d�ޖB����N���E����G��,*:^���=r3ꏚ���d)#zƛ��L˨q�� ��%��m�l�<r<ܛ�߁b�#��Zo����]��Bf���I�jjj��Vu�g-])�Z��ܜe���lZ��ý�J�z�d��l& ��Ti�K�u�_E1;�xC#���R�j��w�唖U mVS_<�e/@@��������ҷt�7�\��r���?Ǜ^���?�Èf}��f͙��~���6��%:Hf�,fHB�Ǜa8L��k�k�V�%U0r�"���f��wL*?��c��y���q����j�������$��F���b�ys`���<����7������&w���s�J�Ll9��̅7��k��cș�ԍ�ݡ�5)�r������ Y���,�ST�tX-��i���O�/#~!!�dV�E�м=����x����pc�`���j���O�F��4��JB�s���;�c���09 ����N�x���6���=j?y������2��T��S������7��B�YL�8DX�q���
� f� ;�{� /���C�\�c�s�2�G{,���T��<���F�.�_d(�p�7=�_���O+����h��R�[�@B��W�)� S�����s� ųT9�Z��C�З;�8���+.�(�wl��K�	��q2"� �������B�r|ϣ"��� �$?Jd˘$ըr��	����5�4��� �m� 1��B�=]���,�/,�������βH��JKE*�.E����{d����ཀ��6�L�ɾ�"-�g��6�khiA}�*�J������Ҟ�@�������>e��nAMN�}�ڬڳ[��F��Y��2'=����1��F��� ۾0v"6�Uxb�T��N�&J1�����_�o����+XF��c܉U��Gf"ؓ��������� ���Ϧd���|�$���	�N8�J=\��oݦ�l)mAGV��C,�.��s�Gd�{��$9�2����H����ȁ�%r���B��ͅ��0��hRV��Q�ࡃ<��g��䇃�	��h};0I�Qc�&v��_O}yG�r��X�DC����#���Ԕ�d����!OO��t��о>M�VY[紋�Q�)�-��]��꫰��y#��,����Hy���f�T�%��ݔ��ߊe2����فn k���M+��谞���>���	h��Ow=�id~t�ӤE��:�.��Ǿ��<?�����u�7e�{�q ={�x� �>�WܥE�>�>��FE�53�.�9��AM�6�5*I�9.��c�o�_�������(�q�ˢ��;���o��ޱ�^e��^/M�/܏��=Xo��~�$0cc����g�\!�4�y��c������_r٭��?A��L�N9ϔ0����Λ��`}?K2\���X�hgxk��.p=��s13���^X�]�������� @�n�����#�j���޴Ăn>g������mck�M�7).��hK�]sk[�-�UQ�2�1��.E�m��̅��Q��S�^3>8ֳn����q�ۄ�f��M�Q@����y��`r�{0�-��@��t�����l��)a��			)Dô�����Ǵ6g 3����X�C��*�
̽[t��V���sB�<�r����v��1�+�e9�m�k�Є@0J���ŭ�<�@�dګ�a�<~ԗ�Go�XD��F��t!�d��-���h�ص5��Ly`��j=}}18�%����BLBG�c��?u4�U�3\@�]b�E��F�����(��8�Ej-����"��]�Y离�bv4M���3G��0mP�q�L�E�z�����բ3���S3��Z���i)�(1	�G�۬V�}�l5�d�6W)/�;g�P{�dy����|����,Y�Ǌ"�S)����ѱx�������bb�����ݥ^-Rm��Ϸ.�����ǋv�k��WQ􊭍6$t���g��|���a��_�e��|�������;U#�\�$}�HX)5ȓD]�Ү��7�ס�[�2�{�E��+tA~/�Z-�*L�M�M�~>��5��ئ��QmG���f�-)�\b y��(�� r�߈3@u�_%[���_���_[�p9_�a+��$�o����t�'|��O�a�3V�0��k
b��d�9�Q!0}�yE���[{GJj_�G��;��M���!͢���3<\zK�龎�z.oy�����]�BcA����A��k����[�Y=̒dL��i���Q�c:��[��k�U�Ua�)�w`w�u���q���)ѷj�j��M���9	���/�!���n�&���~Xf��RS	�T���7N_��L,E?���=������گ��q4�n��<�TߞY�Cx���P�u�zJ��R/��c�^��cz���e�D�|n-���J��;l7v�Q��KZ0*˝���>���w���Q����M�&M_�*2p��<�[�x?�!-�T>��䠀,T��YA��ÌR3�R���qYCj�\�Pp����J���)ϱo8�=��UK���E�go>�G��^U*���CS���=�pN�/}�ɓ��6V�=��?:��R�S�_�7&o���HU�dc�A����[%x6�ХRf�6ﯿ�'W=_9�ܴCD�^����S��,,���q63��F�,�7����FT��J����<JB|K��$v R1�A�'�{��r�r�S���;��MjS��0���i'0>���,�Ş��&bw)%�g}�nG+Т�$&''eII�V��M����[������Pnm���vJ�M
��Ø<�w��s|�2R�g���s�N �ӵӽ<mh�a�ׯ�w1��v:�ͺ��"�-�Z��f��\Q7�1�����3��/w0#����`� ��H�6k���A[/�ډ����|ɏR��d�̊��D��e��"�F%?&��r�Q�ъ�T�kg��q�F���6���ږ��y ,�a�F=�0���f&ŲZ�WPW��Sީ��	3S�G.�$G_8u�<<*0W�Vp��]VvX�7P��㡟�OܵE6�-k@ĆX��E_���MǏ����}k���Xf�W��ҫ'Y�L[��}������a�˒""@��L%��^ ^]���u)IW�ZvVF�=���S.������c�G��^l}tjqS��@��h�w�V���ic��1�#YTH����̝`�iq���b�=�N��H����0�q������VrJ4y��P��1�/�*�זp��jS�B�)����+��O��%�� �cyy�S��F2�q�i��R �����R���>9�:2��qQk��vsh���z9����6־���5#��,��c-b&�U�f��g�(��8c1U�U�����n:PY;'�R	oh����rĄ�H�6��ue�\�$�A�D�����]��e
��h��_�D����20cь�6/�&*r�ݓ���[ʿ��Z�I��c~e8j~��<�X2�=\>�	ί:�:Z��]��/�̸znDԠ<�S��e�#��t��H:32.M�'w�����U�C?"��܊��K8�RZ_�f׺88c�!>��{�Ves�-�r!G
#���5���@>��i1�+�U��A��Ti���fnj�=�F�އ�
��r �l�=hV� TZ�=\p�`�Ac�Y�`-=�y|���x~����܏>qN����������^I�f�H��>L�Ι��P���'�1yI���p��<� �gI��pk^�YZ}�	qj��K�7�`U�K91�1��V�bǆ����N���2�&tS�r��}d��p�ڵ���?�o��ݸ:p�S�ZE���{R�\����cB^0z*-�����_t�l{��b�N��L=����?w2�df��-�ml�Y �fO����p�8.�/���V��~ ��!��VU]#�"�S+i��YD���7y�~L�Wn9����������7(p�Ȕ�.�5s��o��]�(�>V��B��^2�Dz(�M1C,��?FQ���N)��g^��i��kL����p�O�Z�C�kmzo��=gI5x���"=~�S3���mm$�n����AԽ��ӓ}m�����G��FGˉca����k7%�,H��y(�+O��u�<qA&������e����#ZM��{�p6���F�O�"�@��M�{���]#ϣ������mZ�[���O�-��J7vm>oAH-(o	C�2���5�m�{�,�n�"��Tf�8N���j�MS'5���x�����nfbQ����d�r�0�R�z�F��Y��Y��M����O�A�q�N�'նL�?��i%�Ŝr��i��-�=x��Py���\;�����O�p����F�[���[��5���W���iTN3v��6t��de\�M��3%z8w�j�'a6����U���P�����������p�z�%f��O�)2Ϗ5?�`��$������(�*��e�i�f����|$��#N5�ݷ�6 sQb��A��#�m|��s�L.�pԂ~j��aL�}�`�-�D�;��D�P9�^���	�p�S	~��uX���ZQkĻ��iXyx������������2/����c�OO��4�?�hɷM©�/���*`I�n]4�U2��F�������l�z5��a3�BΔ�t�r��"P�~���!��x����#�!���4��[*S���~=��u3ӕ� ���~H��=\�������'�ͯ��Z���R�5�.ГKB5gB���H>�V�����-��]q���?���k�� *W�5�x~�Cd�J����~�祤���e�����؇���[}�[�5�r?
_s��=���%XZY���	ȟ�5���H�Z��֓�Պ�ԁ[���,��Î��|��D����-��;��?�VVφ�7���?�,ܰ3�x�_ .h̡��Ȧ���[$��"3[_kt�-�����E��X ���"�Fv�z�h�`N�|��~��������&�jȀ�&�M�[gl0�q=W|y�.+��ޗRpV�ʀYJR�꼡�뻷Wc�`6���%|wiz���T����h?�X��p���o���OB����>���tD7�\�rQ{;؁:|P�\j7�Q���=a����_��1�+�qi��n͜�bÔ���9����.w�>au ��4iyy<�yw-e�˙����V?��6�r�ϥ��l/S:
n��v&Ѭ����P�k�t��յ��R����gԍ��ߪ�j�|�H�a���4�� ��NԗB��*(Nl��g۳z>N�ˁ˪�W;�`u�9K�W�50i0Hɤ5��c�џ�Mx�?�b�Ә���iǦ�`������]OHIB��|�fb/�d�7�=��;7�xG��5�gҏJ�>����毛X�V�}Uk�t��4�������+��U���H\}�B^�@,��wf�%R�ݷ`kː�����pVu���Җ�U)	y@�
8������o�`�=T��- �皴I��~��Y^pr||���a�����s��x0����t�u�{Ceo{$�2TA�wq�R�p	��������'EK^���,����w~EU��y�:�yf�h��"S���Q��D���� c9�0��2�\������J��c`XP�u	��1`��J��X�@d_� D���&�X
ph#$��!�$;����f��b�03��B�vI�aR�p<�tg�ZX8���ҟxO�7�~�*o�ԭ�ى�А�#S��K���i0�#�-�l�d�z�ޣg/߫+����q��n�c�����"��~�JP��0��ȗ���"��0W��i��V? $��a�8���m`�W�����X����.%vg3?-]A8M�r�����<�.[�B� �]6�5xz溢���B�$A�}������t�&��?�^^$�g�2�D��kb���ZohT1���/��ӻ/K�h����w|0K�RHR�jm=�x��;�qW����ـ�u�������^�	���м����C�80���~�����/n*��u��,�(_� �̰��U��?I�3rrb�:3h�<ڤ͔T���I����QZ��4�k�7C�w�����u'�A����y,2��	�~�4�y��R/�Ƕ��s�'��.Ȧޛ��S|��}��&v��,,\����Qo�G-��3�nј{;|���D��'����Iؾ�3��H�Z{���Xm���i�?g��߄��p�ۊH��%#�+I��e`�*���W�ju�ݼ�?A����m'�\��lu;�F���N��Ŋ� E��O�Y���ƫ�ֳ nt��w ���D!-��Έ�O�@��YqB܂+j �=Sz�Ѵ#������$��]�Y~�{��
���$��q�D��;�82�s�QU�!]Z4�d�J8iR�Byj�
�i$��q%1Pܩ���>I�X������z���;:2rq���������r4G�#S ˲*�̤����CYY=�g~o���
+�q�{�I_��3����||W��J�B����2;p_^8�����:t`�P{e3 qK;O�O���R!���[F��𞡑zyC@��Z�>EJ���VC����^4�أ$�??#\�����I7$�v��WͲh���~��>���Tv[\�AR�%��V_ͼ�mcW��y��p >=mg�e�CM<y�,y��#�����͈��9n�I�����3��V�YVj��X�$$~b16yl��vEη]��ل���B;ښ)�R~�ѧ�"��x�^p�/J��==A
)�ʾ�Z�H����t o��T-����N��l@�b��i C)Z�ɡ17u&��'Z�a�=h�g��;
�dЋ�״�L�Ȝ��\�æ�J��T�Hw;X���@6p�n����x��m-�`�""�"�|֥M55�� %��׈S=���T��ʐWP�Fl�^�vzS%��(��"	3�s��w���zm�i+�3�2~�\)�\��k��y0lD_�+�E_Ѷ�ɷ_���x��h����AID��DoA�A"]tF��;a�Htщ�w����a��!F��|�kY��S�g����Ϲ�� ��.�S+6��xA�F���@�d�(f��Y�J��5�0q[�;젗�H�7	�2�ɜ��a�C��q�fi���_��h(��yxB<Y�¡�vQ�����v*;�A�Nz��OB���Q��]  �h�r$e��+t-t�@xmk�h&���:����V�wc}�TQ�I�햳ᾃ$2Q;/<|t��h��wuX�s�O�M�Ij2(]���
8��:���]����X�(I��Ә`7�ˣT�վ542:B�s7�"��(_fx4薔"�����ϗ�F6O�~?�ET��~K"K++a�]!J=�r4���Aq�^�8����O��*/_�fd��&��`��rm5 p��Pᶞ���W4覚cJ���h�G�Rڋ9_�4!5�$t��j����S���?�,�����0��фyX�em�jb2b��Ĵ�����"�r	b� �D���e���t�����I#�%%��~X Gg��+N�n��o��7f������)�׏F�_8��~Vm�i5�cؙ]$�;��\攻�+���/�.ܧ˜��w=D� �1R/��_Į��^��T��x��K�q�݉�o����{�'2/���G�3�WP�r�R�}#oo3���}N�XWW&0��V���l3*X��>e�+U�B�͚��B�j	�]h����x2!�2���(���f�Y��H9m'�)�Z5��K)0�n4�Pھ_K�����FYl�V�*��T��"7!�v���HS��!�^�式�W�ѿ�[�#��O���`�	nE�z��'(�.ȵaKHѦ���$6���r�w��󛚻��s+X���+�#u�-/���l��>����}�X�Z���^΢�bH���萆�!bW��F����9&m��+��:"LвFY�QlM�L�}��[�u����Ȭ�j�-���P�yte�;a��b�|MS�v�ĕ�OK��J�p2E a	w���9|޷`����n�6U��݇G��IKx�d� ��:Q���f<�����Խ�;FW�\���mο�v�g�����?��g��k���/�U��|C.��,��[��FȺ��U�X%���qcie�͙Wk�����2))xC��
��d�ūv�~�l}�jc����. �.��n�����h?���ܺx��Q!�ǔhV*��!e�Y�L:@�jW����WGC`��U��@s�zsn�{�f�a����WM�����<�7�#�N���Jw���s�;��z��O.�%s#��<1-c�$aq]ݤ۽������I�vL���b����u��s v�Ŭ:fv��f'�C���ϼ��Y���:4�ɻ8�w֎�r�+�ט��4 6�,tA�K_9n9�;�H���;�@��݇�ɻ���0:�a-|j��ug.xi��=��F-^S�n�Ӟ��-I�BA7��ۯ� �X��i�V[�G%�j�&��fD�l�A��V.��}o��5AC�"&/������;ߞ�(gq�I�_�����`*��/P|�����"� �k흃��;���/X�E?p��#]O;�&DRW�6�+�v��|��Q�F�0��G�i�;�MR�5m��D`4�/*�+m@��zs�j ���:�Y���q�	x��/�{�������"0�\����D��������qt���� �����o���ύ��^282�!�`ɣ��ɬ�c��֮x�Y���������DU��� ��g�{�
j�)�#��F�[՛�'[���O����x�Р����
��-�G)(/1͆z�9�xu���in��b��e=�Ґ͜�mh�������G;���H��z:��]��spp];<���\���\�Wh��j���z�;4����$msD��.<�~�!.t�?����7_�&z����p{(�ܨXrн3-/��]�o�Ɖ��.�'dp�~uQ㥺�=-�lZD�lJ���u��ڮ{x��V����d�c�X������oD���@S�/+�@"�z^�%�sh��Z�b0��t�y�����kp
·��X�����&3
ͨ$Z�^-�u�O��Nz�{L<�a*�n��P���nAW�����m�Mr�h	���Yp�?�e�\:�.Os�{}�7S=��_��nib�Ǩ¾xDO2�W�9���S��De0��\�ɴ{��x3�����xn�PD��Ec�+e�"����=:6F�Ζ�a.e��3ߌ><;󬟴�2
���spFn�����y|�:������$�m΃+���Q��H^��[�Q9�$Z�$�
�V!.�3<�\���v?0����Ӯ�
�v �e�%j���<��K���2'U�*��:Ga$�h S�M�Կ�*��ޣ�#�JL�2����X�8���¦�ϝ�bqI���Q��M4i	kO�Ȥӷ#�����f�d�$�k�
H)�������m�[��}�"�-��n7V0P��+���V���6�d�����.�F⦟�F<��}}������7����:p���My-v`7��L%��*�m�6m��｡��?5��<7�#���;#K�H����(S鯰�@�s5Y�g|�c��1�.um������|�e&���'�!�/�3-��<���&
��t0����r�b�l7w��$Vʢ6��6��:��K+e�>��M]]l���?�UL(���BS��W���b��I�O�s�9��<�w�����~پ�	�=�DCU����.ưձ�y��pzһ�i�[6:��+�v~zz��Y7��n���s��vKn��ʩΖx��K_\��7����=٫�a��?�PLQ3Wt�
�?rQ���(Z�%�k6���rD�θ=ўA��b(��T��w\��ܝ�96~�O�_��ַ�X��m�%�hb�*�&��.i3&�$�N�3	�5����f`7��P,��ʍx�}Q�4Q�%Ϥ�'�;���͂�2%s���t��e�0���'�oF�+�f���q�y�ݞx����(J�����o�V����'�~����[t�����	d��n~�U;Xۍd������y��5���*5�䇑����5o<e�zQ�(�Vm�f��ߐ�!|���^ F�Ve�e����?JT�~kϻ���{��Ǯ��7A�
9�n��//F2p�c���qc��}�A�b?�?���z�* ������s�c�)H��`�䰾/�ᖭ��sjx���&@����E	���e�p����f&���^��Y�����uG�J�-	��*`�b(��dk�gs]�aa�g&f���+���Y��=/򁥥_�w5��Wv?^��x��ջ���#x���6B�.�G�'�3��R�IN���b��Iڦ��g���[�ȗ)>U��<c�8�8��׾=�'p,��ۭ��6+D�II�l�*�{���WB�Q�d�Rw�nK9t.����)׌N��g.l�>�;̽vs�ծ,���I**u%�U�_�g�a����ޙc>�k٩�4���*��wb�C��l�@�(��T;���$������Bo[�s���hh��_K,�J��D'7{��fc��b���h&xx�v�k㝎B@��r��F��)6�r�5�&�����?��(�R�D��4�d�]�h�-��ֻn��+���s].�;��6���[l��l�a�?�n��uv�r�3�4���<������G��!Z>Y���/XI	~�z���ʵ`�S�����R6F��6�[���BJm~ｷc������}Im;R}Љ��t�x��7~x�O�v$=󷩬*���wJQQ��=��EW���OR�ӻ��J����x�l���eC�F���ވ���B���_�.�`r�5��?���U�z��H����:�K���ξ�¹����1�D�>��8-�,X�z����Gm�t��QTV#?�7�otS��B���F�xg��[�$�+ ��D��{-�1�)B1��������ikf��q�ߙ����Uy̷���>�U�I9��?�(`�����P�:����n�����9w]>w���/\�%�}W�=�&˱5>-�81��?IxC Q���ӪIm�Ē����9�B����$��;셖^u����󟓵���V[m��d{�	b�֡�B�'Ǵ�]�������¶Ɣ!/.GOoNF����,��̭��v۩@���u��V�0�3�п
��g(9��c�b����5|�����=;�!""�-��lt3�u�aQI�n�M�}���B���e��<b�M@�i��F-m�eZ��J[�c���w������^����{���Mm@�����O����}��S�]?�ĵ�P䟃<ͩyk�9�M��$Qځ��v/��-v׺ןNG��q�MRG(�H��wp���҉]]��[�.w�2���,?���*��[�罳�)� .�a��2��<�	�e�I\�����^)��@
\���(�<��>	��\^X��������E��3z��|��g�	�N�$�h�<.�f��{�h�0�*H��\[�D8c�͎M�׵+��]��b��� *C��Lbʸ	�����g\FHU����}Z'p˺�tЄv{N'ß+��;�����	m������Q����	3��f^%p���-�H|Q� �=磮[���y�r�Я��E �ĝ�c�.�[��{���[�f(���BjB�0���_4�ƺn�����3���s�i��έCI$�=o
%K��/��ll2�󞪧ر�J ��/�[����:���YI:��^n���m�(�7dK(��%�c-�4�	Uƍ�=o�nǿzd��L/6���&#J�[��&*���k�̫�����|E��Q���S")c��6.�	և������Ͽܱ�<%ls<�*h
_/�}����DWo�c�w �����c��:܏S�����}�MH�+��)�-��4��f���a����z���ի����'�٠�����������}%�����Z¢�=�Tdk����	�$�r��4�#u�^Os:�����r�m��ČC�딐�;������򾠒�v�ۗ�mr���tL3x����R����3�Phr�m�ؙPS��W�����d'��T�+O���ო�#�_u��Sl��r�Q��_;�q�Vu�_�#���/�'��Ǒɨ�_RǎB��Q��m�����:��5mf"��^yEn������Y?L�Q?��`.�ugJ��gW�g��{��]`>�d��!S�	��t�Xe�^bw�b������m6[�"~�cN_�O�+����K��^(���r��7��zr��g&g1�/o�\H6O�$������H����o���nض��_(t|�zg�e�o�h��b���|.BC������Ԝ=���%㿐�o]���OQv���-
Si+=6,���YWR�^��}�;Ӏ����������Cx��O��U�j�\��1��֘�����#��=\�p�G�ʿ_K�wݧ��	56�B�s��l�b[��_|��^9��7�>�|���z��A��<���	����XaW-��:�Rs.���˰�|�����q��J|f�]�SZ=,4����AWJ�m\3����
� M������$�G�V�!P�<Z�ʠo�0�V��	�d��׿;����n�Y������(Q7��] ��n�k����#D�N����N_�W�6�x�0��H}�0�-���#�G�����np�z�9[p�<��%]ԾA*��vY_�ިՔ�L�� ��C
��g�������x�d{��h^�����12<fز��f}q�g�a�3>X����`I����7�"v��aXo���_�#�r��b����;8-փ�p�&���wSG/��Yݮ雫�<c����7v�֞���/��{b8�`�r=��]w.]ݎ�򎝩R�^����Hѥ`����@T���@�o/{,p���~��:=��L��(gM�{0i��s�P������8�/54 ݈��`�G9�N�g�����R��8ILGl��w���%y�7QWgv[l��څ��@�`��3�c�1ݏ=Xsv7#L i{1��Q�F�S�0�Ŷ�/���h~#��o�-? ��*���4��X�8�o�W c�v�8?+��A�T?�	T��1�d�n��1Os.EK�����h�U�|�@��~�����,��d��K����;C=�٘ȟ ���SR��c�ӁPV�,<�{{�Sdb4���<��:z��ΚH�Wr�
���B:SFK��};2�����WM�р�u2�	kk�|@x$�����'��ǡ-5Y&�SZ�d�7Nmc�Wz�,��w�k�bb���;e\�.�?�'���C��>�L�����K�R�i���&��a�O���x�{:�\/����M
�,��}L�z��Ltr����}<ӆ��������R��¦��@�~���v�-�+��j]��QHĳ��	3qv|��_�..:�/$��;�Y��Ӻ�y]l�^�5�Dc&��~!�!�����3.Ŗ���V̈i�����aY��2�(�:q�ήٹ��¤���7�.@�1��ᗳh��[H>���I��c�W-ZGA��s��!�b5"�1x�����U1f�wSٸp����1Dc�{�OMШ�	��m����͜��p�Œ?kῃ�ce�H&Ϫ8パP�}��w��i����G�N<��7�u��e�iL�~m_߭���i�A=.�%�	ϑb�k������Th��+���fGQP<` ٛ�i9ϙ0:��m$3�fgf�П�HU�~�;�ҋNyew�]^6�8տeS1�3p^?8w���*�Ha�~�}�t�ɾ1��O�Yj�����H��!��£�G��E�J�2�\CQ23H�^�ռ����pg}��Y�@*s�ߖ��K`�~!s;+�� �4o�������	i�R/��O�L��|�4�]P�s�ȳ_���ho��C9剽�����Ub� �J�/H�L�g��}O��5�?�^D���o��$�f��)B�S+�>y��.K��� �d}��	t8!�����[� ��֟�8�қ�؋�"�V�k5j!e��"��w���
߲I/��֚�iZeb~��S"/X�V�^@?�����xA��Z|G,�崙ů_.d��ё�Ml?4�g������T�Oug�k4T�MŠ;�KP�,_��f���|6&%�fBh��Y�\��O_-�,%��,{틍�ev<�2�"��;�'q��];�#�m��M���,\d��%�+���@M����k������QS��l�V��;YO{B��+��G3Z�pާ�e�<�(�>��z�@p>�o��ȡM�;�9�h��n�F�%ƀ9��T`���m�X�p�b'��^�-.~�c�P�H�Џ!�Di�7j�#���/]�1����ɽn�p��&`�G�l���'����8g�Ee�!��i������X���ۣo�~OWVzQ�d�-ԛ�h{��3�
X���.w��Zb4�Ţ�����5r����*,aɥq<�
���b�c�=�Qa �'�f��.N�V�
���aM��Ҹ��*�+���[��ma��'����i�@Wq�,ػ0�i�+����)���|�>�G��j�%��pS��@�TpՁW?v��� ��.[�D���vk�+��/%��t(P�!r�l=��Y,T�VW:��0�"=z^r����0An��I0��Zi;����tw�a?ExT"��Pj��g�<��,�jQ��ĤCI�����5���.�����R��	��UV%�L?PZ����4O3��w}#NL�����[�'�B?LѮ�EH؞p��|AmS��څرn��(�������1�Ӝ`q���6��]�O�fw.�L����^sƏ�'z�����}��뢰^9%��~�J�ߦ�ԟ��9��(���0����*�m����}�ӯ�7AuD_�䏞?o�^WW��L�9.T���Ƅ�����
�9H����Go�\�wj�5^Ur\�#�۪���G�n%�iOI�����8 $�
SH��}z/�V��k�wf� z�۾c�"��m+�����F�no�����Dd�K�,tW�e�w�>%��ݍ���߄����O��h�-�������P&���J4k.*�9�-�F!e"��!�<��<4!x���yOD ��������[�6@��x�8�H�Ϊ�䤧��MGiv^�|��õ�O_0AP�$�.�XC��
�/��hz6�� ��d�iJF��
����#�mh��9��۟ñ��Ҟؙ��H���k�H����j\�}W�/$�¿`�
V[�J��&u���7&s��ƞw�h�q����n�e�l�ky�8�n���� �-p������1����(Q?��*�ޘ۶�k}6���'����^�E/SG�5r��,�%�gx�V
�l���I��*��X=ѻ���1~��RI����++�a�T����NiG�3|���Փs�
Ā�Cl���}�9��(�L��E	��_�����%��\��Q�;G%��p�r�7"He�˳"���=����υ���OTr�w�R,qݒ̗k�حO�k�tG!����]X�:f���M{r' � � l�U�ʲ��-�+�?A�cH�y~v��� 1�޳��M������-��|���R���o��@�R��0 ��/I�Z^�E����亹��$��C�����|���K7㭏�j/�ǯ+��ٻ���t��� #��m����K���F��CX��6������2�}R���nm�q�g>�����h||���Zq5Œҭb��te�j�:~�jn������������"�m�d+���
�����w��k;�d��WQj�'����.%ɲ7V�X��W:6x�>M�Z8�g:���ū>�6%�&���6�����,�P�.�4⭉5DL���8�L/j���ө����Lx���hi��X�	���~��������|�GLf|�%X8u�{��,�2d�_���\�h��`x]�;�	X2"p�
vi�usݡ�R|�ͤ�Y�3_-�v�|�F�zW��Ơ�q�؝ܚX�}��J�El���N9|蚚;8��v�����@"��%X4�ܯ6���""�}�=�hΏ���y}�ɱDvo��y����6���h��>o=?I#J���OY2n
|�t��΁��s����o��Q��Oka�Q�/%g�8�����_t����O�����K�ͯ�w����{*_1���*Jm7��o7ѥc��R������R��σ߳�3Vn"l&���϶�&�o�h����]�� �ց��ٗ�FN�t��r�]!����-��jk3��ԻO�M"0i[��-�~9D�Eʹ�f\�s5��]��γ���۟''��+|��-�}�������q�HH�5�����-�ʹܒ��3�� ;:�Q��ǌF`�)���ʀ�3/�!�R$����&�:���+��c���}���Y$�>������ؤ���:I��ϣ�4 ��;��[�s�gζk���$� et/|�zR�#��ƴ�kݵH{n��d��� ���lC+ۧO��g�
�G��A[3���ӷ��.1;�
6�s��1���� 	O���T^��5����|�ԯik�����I��6��<ڐ����T�s�Ο���0R���T��\W�J#���Q��_�aV-�8�$��w��o��X�w��Ҙ\y{6�KQ�@�r�FER㴜h�5��t����o�wZ�����0�o��L�d��ll\����z*�)��uх�p�gG�Q&*�nDH����Z�.f�ݬ���B��w���qR\4��:Ix�;-ū��9��@��������<\'����Bh/ ���SK,Óq9��5 �J-��=�����f,���Fg�L�Dl��Y8@� �����;i8B��0 ��@�ࠕ�"QY�t���7s/ġ(��Rb�i�Q ��!WsnЗj�kw&��/�0ë�����P�\Z_� OF�mL�]�M�h�q�@Oy�jP4/0��j��g<���w����g �]�1|==�\�JKb|`�0X�]��-����I�=���i$	�9��P*aV8���7�F3H���*\���>��aYa�'	6?��A[6лb�m����7�־�#��7<2L��Q��9镫pT�&G9�2���|�Wu��y0�A�g8�*��M5��a��(���u��"sJ�Q�_{���[fӱP�(���ΠMCC����C��;�A��(Sc��Er�*4�F6��M ����X�;��x(�'f�7P����:9N��iz\TԷ!�x=Y�3��}� azD(� A�j/���=s�Ns���fw���l��,R�n�]��������Ŝ��z�����*�u�덟�"�_pmL����!���Xm�>�"v��&*A�^P����ט��tDK�2�ZD>-ٟ���8�AN����q.�i��pV���ǟ�
�4���7���6����o5�afx�$E��M�u�Հ����b}��K��շ�_v���K�v�|T�ʮ~�7�wO�~|�K���H��(@@�W�u��Z��L�^V.V���C,�J�dk������~:`�Jk�m���x��w��8��@a�w�%H�wQ�����t�$�M��W+�RZT�T�>�:?����}��������X/�8��mV7F�%f����n��k�w�b>p��)��7���*4��������9��l�)M�+ޘ���@��7V�$<�8�9e����W��N���yU���'�`��r��0,!�{;�ߺ���.�0���|;Ls�I2mǠ���w��>�\��f:_ ����ʒs�GCN�MӒ Ч����OW��K�H��ޔ��lr�Y]s�t^i��B��n�#"�(�G�yJ�aݷGuì��EZ���UG�
�i���}v'���M����	�?�XMS�1j��x�'�����XK��Mi����Џ$���Ȅ�����'�k>
�-9��b�oB��G�]�yj������l�/�ޞ��`��w|^�]:�!�P�{���0]��i�asU�\�d�D���b/�9ƾah��b�y������@��*N}���{��~#��Q6���s��cL�λ���eYOc�\;�U>Ij�t����8E`�\/��B�2 �����\cL�Dџ.+Ӕk��:A$3rI\r~��
��N8�؈5S'\a�]uO�uu��L.�e�pЮMS���k-`9�,���o��TcY��ʏ�w]b�����4����)&��Z=���K�Oمm4�T�6_5���5]�;�6j�`��LPS�Wv/����*u(��6��ܒ�	�;���&
�lW
��v����@����9�&x��m��kJ�X��̕�1�_��%�i��.FT���Y��������<B��k�u�,���ۺ��0������C���_���3b~���}Y	c�m{��i8?�8�(T̝~9E��h�?s(-�Z ���R�1���ꨔZd`�����CJk��pN�ˣc�"X��D�zU��_�5?~'J�t  U|d�b���|mH���$\��Nҹs�܆�k�_�a*��:L�����,�/wRQNKn��Vy]�oK@����h���i�=4�h}�ߞ㘿�TXxw�e^_W).�΍�݆�[ѥ����a��@��/�|(C0��7�0��[Du���w/	ߚe�9�����"#O�:��rt�(5#�p�����3N1޷'9�v���X�-u���Ru�����:p�L@�R�Шצ�P�=&=�z߫����iAZ���h;�?9���s{#���˜����#�ܗd�ئ�E0���N�m�>�t9�x������%����6���ח|����|�@$�2D��+S�s�5"5�y{�Հ}���0�O���0?5Ӌw�QT�7A��7T�<m[s�`��p�$��7[c3�v)c�S�Ce�[#����R��2�o�ă�f���܂6��l��D�I/������М��	,P�ڜ���G��S���Mgȩ$K����Z6��9r���l��&(o������&2��� :� |d�hR��u��g�NA#Q�8�<yy]P���5z����I���[��ZOJ��Bivl�;~c��#����?5��3�6��]�XY~�!��я�Nr�5���3�^ܻ EP �h�V�O���Xa�v�R�i�
���fy�o���D�W�E>��N�$٬
�Sd#�X�=��Y���S��0[s��l�,K�9Ē�:��#	.�KSzZ�޾ͳl"4Z4��I�7>f�{�r�>)��t�}�\��:='c]K;�4:���������ᛥq�J������2UsQ̛�����O!Z
��2�Rf�߲��&�&[5ޑ�&b��伨R��ąm��� ���T�����x��5��j-:zc���3���I$_�i`�X!��,"�[6Sj4�+�W��CS?��=���Gg���!��ӥ��\y�����.�M��=,d�T�
0���`f뻶������=laUZ������*��z�I^J]퉪�էj���+�X�TH5�Zؔ������0��k�ScR#�6?������|O��.3 jA}w	�*���~�7��텶�~��]&j�{��`��I*m��@�B2��J��ss�V�d��VtmV���ɚk��ǊI-��b�F���xαݤ�'�,+��ь���&�c��t�8[lO�(�:1Vp7g/օ���B���:l+�т��#�W��kt���Z����ǔ^��bI��Y�����N��wv{�a�z����K����s����~9G|Rl�}?pb���WG�9.�^��#��&wM5o��;(0�T�3���ϊ��'���G�6�-d��8?x]�d�2C#�n��d��Ǚ�,<*s�7/2�ʭJ�8�������6�/��V��r�K5Ib�$%$��GJ���d�Y�4ٵ�h<wЮ?��ϟ~�N�	��Lp���'�tpq�)�Z�@qhV��Y39��	�C=�;�fk��U<�f��'�����@�Q"�R!	fa4=|�y$�������R���X=#��  A�s�����v6;��O�P{�6��i��:G)߈�ťj'P2����Y���n�R��	����� ���2��D�V�E���d�BG����@p��Ѕg<�ho��e#�4 �@�M�'Z���ǪvZ{z:�Z\u����72v��������� n��D��K�8:�ނ��z!��?e����i�$�&
U�.�G$oő��$�#
kɘ�o��JkH��qL]��v��C���u������iʘc��m�#��h{����1�3i���6|S��}�,��7�Z�h�Y|�����l�y�D�[D�|�m� �!%�"7�Be8lմL���t/��3��ϱIDX�E�6�E
�2	SrhW�f����~S�ګ� !����E�.��$��xr�����I��
�He� f\#KQ�}�#}g�]*�~z���G����3<�L뚒l��x,�Jڒx����N�f�'t�vޅ�y��Ɔ{��^�`e�iJ}�9�I�s�|~W矺Nm	��ߟ!|�����/����޽[����8�#Ю�t�n�.p� d+�n��A�.Ou��L�ݠ��5dcR�'�mS��㙄�2�d��%F���S��@�U��X�,��D�7p4z�~���{e�C�HG�Y���R���YJcd�a$=�j8������L�h�����Z����d���3�ND�A:�����"؜vg4�MPq�h�幩�H���v���7�P�x�>��g�Y�U[G꒦�q
c�2�����8���Bp�g�`�DiG��	��FT��ܭ��T�����'���i�\�{� 3������EB���F|�z�.@M�#U��*�A�aS��^]5ӗ���&��������Mll����Jˤ�vR�,�ڑ�]V�3��SlO ���,Y������~h!#c�¥@@�v��Z�L.�H����e>O0�g���!��B���wߖ��2�WU���/��/z���*iu�F�e�j�v��������KC�D�*�1���bqhIVhq�?@_��ڬ����Ӣ8���)7�~|�>�O=	���H'�6��e��N@�K�?�#�J<G��_���D��N�@�s���~liMm`<���~��I�T���[?���3�O8�������bxb��*��M��~~�d�2@���(@�N�m� �;�f���BGOI4)A,���Fq��k�ҟԍ��T�#���b�Ɇ���R1Y<��W=&�pP�d�P�����b#����� �$����*�D3��(=Q*�\_:�Be�ȧ����E�x���^?z�n��\�iF�}�85����J��p�Tx���5�A��sV���
'Sp�6��u�뼃զ���"�Y���!�[������im���50�aP��büx�&�yǼpM[��,y�-�� �m��钞mY�Շ��GӨj%�F���"����&�g��	?ݟ�}Aq��lbŴ��<AY[(Fm"F�>k�C����Q��9��D'�-�!�)�;��q��`� ��`����-!y��c�Q�W5�6O���E5�>=�s:���/�.�TX�ƚk��Kμ<��1{��>N"�f)6�(���(�.� �-�7+�P8i����֦��?�I��͉ԣ������J;] ��r^���]x�$c����5�aVL0I&�`����O�������ZK�3����R��t���e "Q�G4��4?�+�Ϳ`-�LUU�h�*�2u�Z�t�_Qջ�rFB���*P��~ �(�N_�b�$��J�tq:czyj�nS������s��iaR�ď��~�w�4�Ѷ|3�^Fd�}P��G���j�L�һwf ;��&3��D�>11q��$
?��L��<}���R[S�[1t�c�)�t?�h��x��ċ(C4_�¬/@�v��V���ǟ�\m�#�
�?�i&鵛j�/�p��Y�<ڐ�d�2%b�E�c��k:N��&���I=E�?s�y��0���X���+D����`�����i�c�~k�]���ڝ�y5�-��� ���3��D�9g�<�h��oI��髭��}�%�������n�L`���M�N�`k�ɖꉤ�>��(��e�P�PIÂ�c�,��T�:��ao�\Hy'>J�4	��rR��R�^ghz�>�
3���Ǥ�Z���ג�*����5����1Rdo,�N�����tsDhn���l��2���З�U��1����T�v���-��	-(�^����sz�=W���E�i��_�S�l8�8�J5]%�=�]s���Z�/O%Ξ�>Bnf�K�K��	/�\��쁫�v\N
��W���[�֢��WR����̑Z�ԛ��6�^lf����$deE��ĉ욝�ᒊ,/^<�`[8/��������b�*�\	�4��Utx�Y�h ~�7M�,�@����,�ϒ4��S�*:�rX�}��|�������h�����>�
�iw���޾��Y�������V����x���ӟ�y�	3�d��k䣉xt:[�	����?�]S��ZO�\��a��zn��y��`��&�ޝ�o9�?6������z��=�1�q�b"U�\`�ɺ-�Bo1�wf~#
��:գ]����4�A��}-mhe��F�����*�#o�����_�i*��+�N����W��;�#�i���k�v�X.@��������0Y�|�6��П�$�灇�o��#L��,��Vf�)����¨AHba^�Bk ���xvgJ�	�]]D"����^�h�����-�Y������pɃ����[��z�B�t?m4G6�û�ďcl+W���E��$'�������Y�������g������F�No�ӻ�?�5R\�=z�[��a�\���"���Y�q�^���1miU����v��#ɸQ��+%v���peּ�w��J��� �K�����'���a00⁺���fdZ_�k�/'�M-Z�%ɹ�E�I/�4+7}�����~S�S���]�ьB27[43##���}DWg�c�����|�b�b�!U=:�c��k���%5�Kh	��c����`
F������p��J�{O�e�X\�����E_J�)��T����i�x�����B[��{��;zDM_�m$VA�w��Ww&��_��f�y*{q>z�ڡפoۚ�h{��Ŵ�Ҹ������H14�nG�]�>�%$�����7h��d_)�[
��3K�W����		� �޷��[z����ً@�j��E�S8�
��y�� �°��i�����;�L����{�42R��"�k���,�0<4Wo�����/Sn%�%eL�tf"#(�AD�ؗg��L��-zT�y�lc2H�}l�"϶Pc��:bc�;�[�ᳯ�c�������Qk樅!cn��2*�Y5{��ؼ^�N������3���]�rtm�𧺹ts��\�q<=3J��S��d��8���b;�+�4״综)тF6Њ<�<]eX�M^�n�IAiDʥ�����S$��R���U�;��\����E}?�x]�Ϝ�9�)��(�w�ԋ��%"�%���o	����= h�]^yK�~�Ww�|�Hf�д�,�/�A�����d-��*9�j��±�P�M7f��:��F�x@8iMrz�����@3��]ډ_�#�mӭi���]�N�V�JtWTg�
��Ii���/ i�@9mY2ڱ�R�����<!66<�+z�ȧA�=�7o�"��x���I��Qt�H�I�B�k7<~¯\"YX��I`,��*�������DIݮ����EG�x�$M����pK�f��k���ߞ,�LW�&�`���[�gM����������&>j�܃,]���ڲ�a���g突O3��B��4���n؟�j����%�d���x��q�܆x�^C�[���3��>����ğ�ܬ$I ��/�U�&D���b����T������c[/B����1#Ȳ}�����ϑ�v���{��dǺώ�nۃ!��|um㑚�v��)�}Ɖ�{�����j��=�}g�� �}�$6\.%oZ��B���1����$�D��z��4��Q�����y��#,X�bY��Fߎ�-��i�ݭ�r"X����-N��l�e
]|.2��;��'
�{����
��)grmc�v@y����3�Í��n�ʱ������VώI�(ݗ�fn�I�y����|m�z�ޘY�&��M���|?ZG刮� ���b�@�#�Kb��edثg�����p�]1Ӷ�O�%�S*�y���FA�T������_r�f����+(�8�N��GK����X��\g�Ш�b�R�o���b����l���� �T�q�l�Xn�A�d�R~'-�����T&s��=���vvt�S�{c��;dOo�=��?ۓ=pmQ�EwE�H�N�e�����k�gf0�Y��܋��	�+�K�K~Qt������B_Z����4jagF�b��G���XNj�EȄ/,���+eŇ��؆#�"��J�^G��A�h0�uʇ変��W�W'[�o��V����ȍ����I-�\Ȁ -��VS�>%�%��Ci�k����TN�`��|��}Kq��٬XG#�dwY"�U#֫�O@���*~�
='JVt�2�Li>S��m�I���F���Y����.f���Ow4���2�X������S.T�c��	�h��9�v���(��o�N�Gxԉ`Q�`�C�v�$ZH-f�<˰� �t�
d�]'{&�`\��ʉ.�ڨo|����,$�=� +˃������X�Ǫ����e�����ė��gG*y��+��&4��v]5�����-s���jx�R�â��M�]�c������S5���%�D�u݀��`��R8�Ԅ�ꪖ��.NqY��=�6>0v��
�}��ހ|O���hJ�{k���^��g���3����(�T�sK7yssé�(�&T���?�yӰɧ��U��]�gض�.zfp�E^l�]K~[�S�r�i�hT�s��h-�e�l=�e�<�ˁ"��p��>i�B��\�����l�����)	&f��g`X�!~��4�ݗ�ykJ���{����r�KO	���ޅ��o���UEj���0��
,zH�c��r��TWщ�-����X���:�#�v��s��+e�����K����>"�skD���86袟�ި�`�Oǃ�c:�]o��Y^	ћ�}cK��T[�bj�k%�Z;�.>[�0���r����7�Z_�]���s�)n���'E�Zx%��q~%L+>�����%�Xz���������1�ޝ�<.U7>�o<6O�|�S<Ʋ��� 6�� dt�2f��/=D��a%:uo�/����5�ӢD��S	�=���<�����b-��[X2�t{RV�i'(�ɮ��q�d�Y�т�Ͼ�t�C#��l���{�y>����r�}������c��L��k�Ԅ�G�p�]w��p-��V&&xf�' �pd��LW2c�x^������k���6�mJu���ѽOc�v��zPKeZ�|���}p�RR�R���QTZ��z��^t�8۝ܞ.�~!�����)5�꺯��@��=�3�T�S��{�,{���`�hHN�3���:Fשn@���%�����yҨ2*t)������F�#ҫ���I��<S�"b�r9��y{T�7�a���j�����c���Fcu��^�6\�
z7�"��m;�o���������F�G R�i���	�	@p�͜�!M���p����g���=�ޜ�^�#uEm�bs>t��)lMN�/9	�o�8�~��&rzxx|���<�@��~�e>��+=6-�����
R]?��g��2%��|)^É(�we�ǰ����\�ZIi�
I6V ,�Y�Î�s���zO��$q��x�s���e��P=!�R�VJEmk��wwM�]��m�R�4fF�g� U"�(%BY����G�g��-柸�8�����/4�g�l��%��74��ߴ�ʂ{bK?��ex{�[]��-:�:�5J�xְ�f��zCK��ڿ��X�@=]Va����l3��X ����ѕk���ŉ~(�MƵ1�+����x�=�k��G�+�;� �а�lU�)���7��� p���Q�)�l�
�)Q�Į�`Ӣ-���z����f' ���z�⁏�-��K� #ee���W�b�D�?�@Z���w�����LC�u=�%�n����F�����L?)��Q�-[�|������V�~�|�)�����NO���L�I�6w5xb,#4ǯ�R
��,o����
��&gim��[Bw�����Q,���!�7�.��m���f�P!�"3�g�ig�B��u��o:�(��i7!��Tj���K5�0�??K�3��N�?oW�r�T�Cr��xB��V$���ڵ���>^�x�՘ۋzi[C�d�&��e��yc�p����$�^J��o�����RkI:�����h:�(���=�X?��!�R�i.gvݝ������j�푷����Ҳ?ܖZ7X2T3�^늌���Ķ����˗�?��]��}oM̥B��щ����)�k��ӎ���<�Bz�w#��"{S���&�'�z{�rfI		�yZ���W��[y��{~��EKk:y�a�����b�1%kHFWg��WVl��Ȓ�-��qkt2.S��IMK���Gx�z�.OU�h�!�6P�/�p��͠���K @�:� -}��I8獣p�7��1�[.�|��~n�\"lR9>��(�e|q���fo�ް�Ɍ|'�E�3�i5;Z�nI9�@%@>Uw�� ���O��׎$ͤ1�f��x�>&�@���$��>X[M���`N������|��@a�MOȴBi�մ�nΒ7���d�1,	�8�8���_��r����}�����Y*&+�m9�����0�Ѹ��K~���]Ȥ���.��9U��Ѱ�dj
����?ۋ��W-kQ��u�ֺ�C�Ep�,x�-��Mj����5`�Hs[r�������a�n��Dpu���b���zr�����ARL����Adi�w�۰�ބϩR�����V�\����d��!n�&7��j������Q7���|���5up�zUp
�Ȏ��εj�!M��H���[/�/��9�,j5�����%" Q��~��z��<֌6�3B��5��VES%�J$$?� V��aF#��Ԑ���Q��ൂz�G���,J2���>8u�WOzR���)%���~��d��Y*�ˇ�D�{e�<���>���������8MN��+� ���FW-黽������c�E][��Խ���a����syYe��nn��k���k]�V��9R��j��n�]:FîvA�AO�����i�I��o�z�� d����Y�h5nH��]� �r?۟(͜��Q$|1�HS%��6hI/�0+�<=�P�j�Y�PQF�MN�<���<�Q�ʪR$�L�������4�7��Q�}���?�_�Lj|ob�Vs��w9-��2[��.�tv5G�X)U{��R "N},�Tl�C{�MF������9��p0����k�y�gnʻ�=�q{,zLe�suVK�zc�7���RZҩ �C9�7'���M}eʹ�Q��y.'���&�_azӶIVe��K5V��3����q޷�k}�Vv^�������/����Z������y��BCcD)��Dv��[�nu[�T] �c�(Ѫ�]�v�q����M<�Ϫ��K
�f��%��s��R.Z��s^=����"5O��R܉|�xvv#u��(
;;��_s*�	ڋ蛟:�R�q�ጇ#�c}��
mW�?���6ԯ���5	B����GG��k �.�����C�+����t.~���W-:�Ɍ����RqoN�n��.Ş.��WdE��4L���ZZc��	��9/�y���#B�K�4���f�Z�V�\p�5����y�lL�]�h�M�J̲�����_������n������ZR�m}"f�kD=��o������[	����'�MrY3ؙl�߁���b	|�H�B��M��>v�D�1����/���%���.<��Kޜ=r��i���V~����=�`��d�D@�q��y��c�Vg��ف�~W��w�J3�tf���L/^O�P�,�#�y�"B)�����c�����뢈��B���Tz�Ȼ>��>N���1�,\�s7>����I�.{@f�W�'��Kx�U�n�� �kT�D���̻������.p��ާbi��mQ��y�@�����?�^Q��p}���<���$3_��C����FZ��5`[ӝ.c���UZZರ�W&�3��ew:��Aܔ�`Nw��L'�.��ӝ�Q�h�/3��L�u�?���'p⥤%�e�f��)��'v��{C?8?I������म�Eq9���}�f��6�9.�0�)q�jpH#��3́*h��_��JS���k���uC����|�迳�b���C2�|���!v�����E{&��6�30Q���/w��94��#�5r��7�+>WKZ�s��C(��>g:�껎�P��^�x��|�h��9��B,L��$�~�H��?rZ���^*���DqF9a����ϕY6��ɢb�C�P��ԓTr�{/�׻},�>Ңy���0�Ò��tG]K����9�k@��޶<��7��Oj�{YԀ!���trVk����G�ڍ5nؗZ�[�&����D�V[� -���,���>�}�n����;���<l��ah�c��.�h��߭�q�}���O�.L&{hRͭhл�"�U��?��y+&1~�X�Y����&6T"i�i�C��U	>j?��|؎/���k#Ӌ�RO�02߱��i!��ur�Џn��L�"غ�(H��'K>���+�xZ��7��N3����!��mt��"K��}{\%�->Z���F��a~�*��1�&cl��b�oͥ����ݬSlex���D�ib��4R�6h��DR.�|P�F����_d�J/�)��D����?�����W�bB�'���^���X��)��iN/ZІ<~�nQahGQ�7rk'A�������|DJ�%4����%:�{��z_��]T�Ǚ���y�c�1��d�}(�P�����2�����E��E�X�9����C�*�xl?�f��C�>�/�)<�3C�@nv[0��/U<$�7^W�y�UG���y��4����P=^��v�cL��(�mlы`ܳ�@D����� ┿�(���ٵs�(��+�SaK.-������gNC�{�3?�w���n�ɖ玳�%�g��#P�/�<�F�εS9��&�d�g��R����2�|�hjɅ��q_��<���0�*G#Љ�����'���!е��SHѮ$�	̐�j����;�"JZ�iՠB\���-�]�_�w�S��ӖC3�5˱+��"�h��C��z�ޚ
3��l[��+��oqk`�^Hx�����)RaXn?Gd��5�Ųf��D����`|���[0L�]��R�I�(�7�1�,���װ�VMY�
�f�a�k��'���������o����d���G�3.N&N?K�7�p����6��p./��.��#f4-l3U�+p)7$��-���$I�����C4/�G3�|��u�3z!��Cy ��E��SZ����N�����r2���o�����/�Č�_:�v?U�1���C �lÏ�wg{�? �¢�hyUNR*( ;���_�u/ <�6y����ZX���S)�_�lAa�T:�éڐ����M64JJ"��a�ng.Q��� �ܟ�ؓ�at*��^�+M���|06�tǤ�\�B	��xۦ���H9���S.���؟5�l���H>׻����·(���%��0�0�?���DF�eK"��>��w>�	P\n��0J��;:��`1�?(�I\���b�=V�Q��j�y[gh�NX��U)v?�`��{G1a����Y��B��^��,]ng�}���L��JGVR��-}ಙim��*�s� )M?�&Y�n��ؙ���p��#  '����bY�B��n���O�"����罫�B�C�Y�5�ڲ�����~Ȭ�[�7�|�$��1�k7�v�Jr����j�}�H�$�;���6��芼��@H�){dt .9po�L/�W@3������ln/�3�9Y[�Ĕ��
"}��*�+��>>��J";3J�}ۿ:�sl���`��gld�w�\s���)[���w��ߍR����Hn���C�,Z��fX�Y(�eT���^�?�,�De뉙�y��*z{�w��\\��nq�Q����Ԏf*���Ѹc9�4%��^����v����#Ǳ��&���Y�=G���qH�+`f�Dj��2j�w^c��S�����=��*�_�P��t�/u}���@ɰ��c�zD�n�ѿ1���{��nu��S>�[���hP�%�F��+�F�]���c�I�#B����b�U�����Oe<�]��n444�o�Ę�K|�DJm
%�VX��+�kf��ghGj�W��E��_��?يu_���c1����ȟ�T
J��-�Z[����~�b��x��5�-й�����F���Dұ]����;�A@���?M����v�c�p�7E�X	�_0�EgsUs��w" ��V����'-��mN*V8e�:��C��rW�|��������_�6sUL�}���e�)pq[�v&[G�;�	�~?1�ڳ�|'W6"xXۆH�X��gX����*�Wo7��FJ@�ő�)�񝚪L~X���Ok~M9�o���R���0DS��}��B�6�'W(P����A��wf*{X7A�qΈ�+�����a+�uM"��.��2~[�����E���Lc0���9�PhG;��]K̈b|�&��j?-O)�����O���5�Wh$�+E- R��˿���W(���WN{��|�Q*�*���Ͷ�>:�~j54�W�L���i
3`}�m�%�Md�`v�<�ߢ��Hli���Z<*��3��|��jB��@����-��s��/�>,|�Q*��RGS�`$����ʤ�U�7� �Ė���������1���!��u��d[BOO_�����um��ˇ9YL|�XP	��WZѼ3�_y��EF�+@���J�a	M��э�����~�?R��lі��ʶ��Q=o"Fҿ0-E~���0+���O�����g��JW˵�w[m����Kӌ���KE��c�BW^���J�D�,X���?ޜ��\� پR��@1)�q�fyyq���-J-N�L�A�����kn��A�#����W���^�9%߾�j�\����zq�=	��\4��B�ۿ�S:�!Ӣ�F��{F:��V0��3�P����cR����\d^��"rD�3�/j�^���,26 �\�O�G#����3Yp�ehπ��sX�W�7�t�K,{�f)]e�z������%�n�dg���B����v�h��x�}�+����[t��}5s�{��$Ð�����ML{3�G��_���{�����s��W�l���ϊL'��f�0��l�b�)C������J�ѻ�c[��d#:�zFF��a��R?�͵ܖiXY�`bd<^����/~��)���>%�O�KWZ�W߻���:�3S	���E��5Djr*�4�^��: xk\z�e�w��tK+P3[�b:bU�*y�HN�S���S�4+��&��%���8����B�����3��4�9Y�эVrά�h|�{��3������+&)ޛ��$40ee�I���l��-kܻ�˄@NXDҨ���O�ާ�u��-�C�kq�/�/ r������Zd���	�Q��>ed5�g(k��̧aϑ:hI���?�Lr{�w�E�+d� W��A���w�-��_}6N4�DE���5���k������V��|%r-sY�*��ޗA(xr��.��7�F�(��H����)EU~}��_cd�^�/)-#�#`���\����Ԅ�;g�$(���[*����A^����(XIA�F ��1�Aa�^u���	@��:��1j!ʮ8��s~f�:��p�R_���r+>����Ɯ~rM��+��Q�~�j�$���	�ㅫ�U�S�g|�Ȫ���9`,{s�}^K����`�˶wX2;w.ŧk^+\0|�d��]ŭ'V�i�������F�l�,:�������v?���_���o�����M��ڑ1������:�����?�#���4J�?3�ͼ$�����&r.>��'��e\�GSZR�TÀp>|�9������fF�Ɏ��+M�Y��K�JKZ�F�B���ﺙ P*�קKwW7+�?&�Ve*\�)�b����%3�5/go�߹>��j�ӑꗊU/󢄼�-Q��L����R�J��Z���8p̘�>ǃ�9Or=��|c����E�r5W*�[��e��)�~��K�N�-�����~֐��w�fs�Ҿ1���,���ΘH�+ئi�)�i��<�	<Sqs`��p��e�_<ܟK?��ɿ�"(�S�cل�h�MھNo3
��� �ƦJbc����=(�ޒ���H^D�����5�+B�q��O�DK�C��<C�j1���,�J�!K��I�#	�G8S���Hty�e�%ى���)G��鹆�"��H��"��a��R�w�-|ok�� P���^��qR�]�T���[&Q"�E� �*@�W��A����фh�.�Q���w��A�.�G<EU-f}w�1���.GSZ��7Ԋ@8u�)�E&Kq��AZT�>�����7�D/��S_M�{Cbu�������E!P����/���uVy�Z7�dQ��Əz>�u��6�; ��#�ù.��{���	y`��9�t�.X�E�C�L�h~��Sc�	�
3`���즿���izH
�� ��`$�h���K���F5@AO�������ϵ�k6�_��4ʋ�H�Ee��_
`S!݊96R����!��M~-��?���`d��|�����]���NᡏlL��P�n1�H����>��c�]��
��-��F��hw��Eo*���n�v��}�+�%X�a��/l��3����i���&D;ykm@g�NRL�&6rW$�P��IV��q�rn�����=͈n	�¯O��e���wf7�=�-a��	��i�uq����W	�^�g�V�U���hǲ���y윚�	b+�	L�އH�v�#5E�מ�w�h���?��nZ�(���Nh5m��~��0�#�k�$�J�AaL�៲�z&z�G�N�t��L��#o��m	�MV���6����J.՗�����Yq���s~�d�,K�v��
�(���� 
x�9,��}��+ǟ��^ ��!)�;�[.���X�p�UǆǕ&D/�C�j�;�#i��hn�O	`.�H�j�"H��$˖��X��ddi��� VZ��X7�s�U"�W�[�"�����Gs�u��[A7[1����Qx	N����_�os�7�,�2|���쇃�@����7.��l[G�R�:��/�	f����Ѫ���ԙg��ؗ`��ܪ�ڼ��k<mj��M4�v��օ���Ϗ�ϓh�W��f�b
	%��"e��ws�/Ϳ> �1���2YW���a�m�!迳 �Y�ѓL�H�J¿3�A��!�Xf�r.2��j������9�����:����m�O�[��4��)����N-��ģF��%�"f�L�V*y�a�7R�	}�i^�.P��|{��4�Y�)�<(�g=Irh��g�B�sWJ��7�zߐ1V��U�ə��9�q��/�61"E�C��*��g�7�0��<�����a!�r旁"iB�[O������q�ߍ��_��iMah���.�2����;�a6��C@g�t���9��k��T�����'�!����g����� �����)_�/2O�{ߎ*�j6ME�r������"}u���&*�ce\�*�L[��6��!�XN��d��m	�!RQ���k����i^�������"Vor�������c���O�j�0�����4���X�na����r�{��s�f}�0ڗ�Gp?;2: ����#/f* p�
s��i�g4���S��[�4��̌K��d���'iP���t���E�y�������@��.{bMd��`<�|M�3�d���#Ӏ������&�o=�.��L�(�@��9'j����J�"�x�&g�2l�%���Z�ZL�w}J� ��K����:;v���;(�_�l�\?�0�}w�^�t�)�33!3d;Ӑ���T�bt��5�*X���a���\}-�8Y����x%S��c�q\aJ�ڀK�V�^ !����� ;*ŶV���ˏQ)�[�Y�B�sG"^΁R�� �w�Z��qM�rf,:~��Ӟ(��
���q
����gcbU��m��o+�X�!i6��?�s���ּ��c��t�!! ��
��
�����s�]�1��Q�;|���V�?�������{��߼�q���2^��mn��G�PF���g�o�+_�� b��GG�!�aς��(�@�B� V�o�C�f%�f"3mK�5_�:Ǚ�y�O�XH2��2��3dI3TL�|vs7W��FVJ���)��\Ї�@3��(.�7�O�Mͦ�b6������AG��1�0c�?"�)r�]�
`�(��k!�<U�گ�qG�Cf�Fh*ڔ&�nN	k����5���T�Q�h<����(��C �4�;�P�p�XY5/c�E
B�C�ە��R>�tC��p ��u���nz7�w{�V���:>	���_�"���沲ȭ�R��=�'��e>�c�s��X��\O�<��t?S3x����ֽy�]�g�%7:�V�̀�k�o�EO��M$!|6d��,�-M[�0�=QJb���A;,<�����5�|r��5��l] �?�SP �JG>hAN�;�؂�\tG~x�b���c�{��@�UW?���?2�!� ���23���C�����`Vѱ��R�%F���P��� �9�Ƈi����7�ٍ�׿����{���H�<HzM}���[�����6�ӓ���[/y�4"Ԭ���}�Ѩa��y��w��� @&>��~P���(����ST>vP��?��!��B�,�4��_��h��h%�N,� R�VJ�psب?��WR&����E�F���T�66�S&�{n+��Ȁ$��%�˿Q��>tG�پTA�ƯB���%��w�W�������Y(���u�7�V�دXd�8~~�Ӻ��O�ҝ���-#�MB���������C՗d�@�~�@�P��otii;�,��хM]�{���k!��Di�k����kt#e������[��1&�#��{��r_:�;a��l��E	b�q��h�B	zMzn+	|�ub�p�{�Δ�]��mI|�����Y*��K����b��\�DX+.;���#2�0���;��Z[E.� .�Ǫ��|g`�Qj��+)��O��a^�	6D*��^L����젻��I.� f[��r���O�����FRg�-�
��)�Hӵ�Y��)�}TH%��"�fuOӵ�DXV��
��Ȅ��8��s���kj{����ǄΕD�U���r���{x�f�1W����lP�Q2�7ih|���? yЯq"_"
%7.�S�!2:p��N8O��#�k������E�J���Q` �h^�L�_t��@�3�����$	KmsTv�3 IM��KK3���Rfk�/�R�v�r��[�vﻜR=�&d����G��v>��B�#ӥZ��p�kq��]������`�e�8�́_�Zt����N�p���`ְ�㫘tv[��-䝝U��$�Zn)�?1ݏ���ZGB��sG�H7#9R���l��z�=�� ������LtBﺋ�������q�{�mk9#Q��q;�Q �k͓?�8�*��x'
�q(�f�|�b~0���X����&��xL[J-��S�sm�����ܟ��u��ў����K�E����	��K�i��n1j���	�����J�H�:Ѷ�����lz�T��w�NM�E,#MP��|��	܌w�.�{fX��dZ|���.��"d�V�jk�x�g�v;;`��\��ӑ��+U��d�H��zQ�H�,G�N��׭:w�ܐ���V{�j�WB�	�:�"ɑ��`Ё�ZƵ��ֹ��f�����Y?9�x�@#H��D��#"���֌-P�7A��PF��g�إ'<���K�_�DtS�%�.��C���B۲7X?�N�uGw�FGQ�/�z��#!\]���_�_��&�?"!a��c����8����&�������V?{�'�}��[�m��X͚���7#qI�}:���(��%�Y���̏M3�ڳʜ��*n��V�|���N�������|j��؄*d���h��+��R�(	����: �B�Ջ�[�7~{2����v���y�-\��7�&�`ZϮ1��}f�g��U�`�ǁ��.L���c�k��8�\���QF���?����>Q!T@*��5�H�IV�B���Պ:b��r;#������i ���g.&�����W�-u����	���۾FX���������&dz�h��E����Ô�	�s7m"Q�O>��Ɯ��JEuhy�wx���y�2�Q����Z��)��:�I&C���o��{�)���*���r!�q����ɼ�S���a�NK>�f��b����/�^be~�:+VW�����l�&8Vm���K��$�a{u�]O������O=r�C ��;��@��������s�����V<��5����y"p��m�����w�@�z��I�@Rɟ�e��ț�x>��Ly��J�\��{�΢���+!�*|$Tlw������w*����\裦��l��|�`��u|���kw>��;�}D�w�ǀ\cE���,�5�՚ǮU-���o��-ٳa����ҭ��E �6o�D�q�t{���������eO7�6��^���J��H�\I�|�/�R���[Y�y
���bx����W�I�9	Η�:3�_�7Z�����#d�[�6���� �ڒ��{�}H-���__G�!�3m���;vS����"d���HcM��W���&�/f�b�/�f���������^zV���v����"�E��b�%�[GF	l�U���nXu[�)��+����[���?.:�������yq[d�������9�+0K�� 8,��ⓝ�I�+vDz��K�\�_>�����HZ�6�@�UûM!��*����GJ���A���$�g����������Z�AV�J����$�kQ���c9vN旫Wr�=9��=���E�k+��G��Yp}Q�DǄ��1�W�H/= ��dɵ����zM��m�nkb���8����So'��j�h�se��}�n�|����0N_�G�eT&���{"��"ƕ��[�)����Do�O���5KUw������(�̖��NB"�37S��[�1=N??d2�떀j�D>%����@y�6����EhI�[%�8+Μ�)�i|\T��T���s��9��%�<��IY���Jq��
J{�VT�;Hw4�7
�͙�Mq#B�A-U5qby�)�*�A��}����Y�S$���l�h�bˤ�5�	�ڹ[��̪�2�J��z���1�R6��;���s狟w�gz��8�<�����J��>8��Q�c�%�W9�j*�@�OA�2���N�0&mF~���n��N��tdb/U�i�<� M����G��8�Sn;4�(�6�ٟr"�T`5��zJ�ߠ����1�4K�^�%��)���墲S���s*�Y�k�Uk�oR`�������T_>�T\���?f������a���j��n�p�b��`B��M).v�YYH0�ʼho.-��zk�pXu�Q�:���74��՟M�tI2�Y�`ߥ$4׿��`���}�v�ʇr�/�Җ���)�e���'�g�� @JI���{�L���f挡Jv�X�`<�(j7��BTR�[�|��m��Ѻ�u�3���$d���}��5}w����Aꛝ:WW��NRx�"��B'�G�ı�$q5�j+��_��@�,��X���A��^"���C��ȃz�{T�~�ߟ`�$�����4��V#2P/S�&��Vt��?�w7��-Th���0 {!LF�=7�V��ؙ��V}�kE�ǥ�"p��j�̶�r��W������r�W��rv�)�Hp��V߆�ߟ��a?8E]Q�dM�X�l<e����F_X�R�K�C>�V�y����W�%5��>�z)Grߢt�$F��q���%�@�~� �S,k��Rg���Ǯ���u�ީ�^'�?9ـz���N[� �`cİ�h;�b��^pC�T�X�+p���%����{p���b�y5��}˧�t�g�uH�����/����ŏ�p~��ʗ����I�����V������^!#�Y�ԪT��g�e�c��<\ؼ�K�b{f32�f�.!a�H/�b�GA� s.O?�:6��=�����4�f��b��L�|&�!�&(L�(+�F}"%1֭�?^��"y���hﱆ�,|O�����7q�0L!��.����H�>�e�����mX�O�3��%��+�VFb��%x����$�W��$�HAcB�n���ÒQ��N}���F!�)-, `�3��!�j���J���˾n��,R��i0l�����{�H��|5ٶ�����A�Wʮ��� ��6���bo�J�CɊ�F�&!� �Տ���3>>�s E�n�Rh���E���I��;zj.4�D�=�9��J׽�7��_T�%�=O2����/�F޺>>)�RIwI�7�d��a.RC��s�,&
+�u���0�֞i�G����:�z���霪��c��h���}N��D�5?2�d�I���R��ZH�Eϣ���iiYd��Og��T)*	��-X$���v�7nDq�bI��-I�a���Fv�����)��{��Qɴ���N��|M�9
1XX��-w勴��&X-��F��Yt]�u����V�k�Jg�Ҁ�{�Lx�3N��~2�|�����]ٶ�E��3z�jl�����@t�|+YBW�b�#r�k8�ᐦ�.]Ȫiw�. M�L�oY��ыm��>M����Y��
��op�R��:՚`3P�ݞ�!w��2������.����/�a���w��G�E��U|cﻅ~R�.48(Fʅ,JHL�TV}�S���O����i</�����-�A���o�k�*KК�z��H��B�c{
c�J�(�acNDK���SO��\�����-�-��K��a�;�6�{��)�"��{i��&T0������"E5+acC���w������6�f,.�cVό7�}_ACt=�]�/��k3�ו�R�OQ ��`}o�>�-�ju�r@���m���k�OP�;zF��u�ci��@���TT���M�Sa}W��\��Ύ+����%�e(��J����O��&%�ܱ�D?4�Yx��U}�O���43�Dfx����fk.��lKڪ}���Gg�����"��}= X���C��Gy�sձ�b���')��ja@��Ѡ�/�v��!�:s�<vS$B���:w\���*\\�ʭ��Z��+CH�����	~'�=΋X�Z0�1^�ٷ��2~|?7Ӥwv��z��U�,�3�z+�|���V
���<��V�>x�Ȩ2�')�.�\��C�rۍ�c�����?6B%�A�m�_X²��p&���U��ދY}��N�]߯z@f���ֵJ:���W|���s�_�,�(?�m����v$h�B�v{.�n�/j�W��8�?������ �:#���2�_n{����g��h-|u���r��rBV~j�!�	a�^�F�m�鷣=�?xыmS߸+^�<(��Ƶ��cL6��B4��2֪�77P��^jYú�gQ{��$R%�$i蘔ޥD��ݪ�~Od]���)Pv<�)\h
�K�	�����鮬���7���"�O|��/�vn�\�������� q��.��_}{��cEwc��tλ8׆Z�b����Q�?������2i���0�Ƅ�
�{��R�*�ʟݙ~*D�}D
���H'��'�5Gk��L7d �7�a"	L�*O�(��r�5�t���|��d��Q
H�-�Cc�?��Y܃�h �V�~6�O��x�A(�mRT_�%|t�������k��%�A��n$��!]ҍt�t�J#HwwKw(]�����;��{�yP;f֬5g��Y�GJe��Y�*]������C����lh��[��8�0�����H�prg��7U���;�C
�r�k�����"$<�5�'��-O��U��:�ϫz>4e�gn�I�M!(���^/����������_��͹������c�U|+��9�W����������B�dD���?2'�gMx�������;{��<�ғ�?���<��\Sݮ9�񗶬�E]ጵ����\�}�ݖ<
����\��\d����o�Q�D�e�����ι��el4h�Զ��rF"Y�v��y��㈍G(�Q�%���3(�:�HY}$�Uqa��,�Z`��,cK���S��4݉�A^�)S� ��M$�� ���[=W4���L_88P�+�����4�n��m�da��x�����f�!|�;˘C�{bA��)������ܒQa�	#)��[Go����䐗��|B��q:qYn޻�-��D`�;��\eP�%���ֹ����)��,�댾'�K�Y�v
Y��[;e��<ᓯ
���XDq����Q����^��/b��1*xx�����~�09C��2cwvwo��@!��YO���gf�dad��PS��do�hwq�m�\�f�ȖJ����5*��	]V��$��Ӌ�>W��R��x���N��r��q��F�4�Sf�yK���G�-�d�}��I�����j����s���	��/�f������&2��~�V����,{-�k�?%9����չ=r�������� GO�����g9Vb���I	ʶ�z�ėڪ�if�C�*^�=�J��L댭�p���~)�U�(8�E?[����V\�Ɍ|Hh�+���W��z��� ��1�n+G>ӗ=���E8��t��~wwW�����Kp{k<��O�$�"@��:�q����@ߍ�NM�E�hx/__`5��L�F?3V.9ǖ���=��N��g�rM��TS�f�wc������3�wr�����c���o*��0^7���٨�xD����x��&/�R)�P�w�ngy�h&����u`��R6ф������4U�0���q�6�PK�h��<��|J�f�L�\���a/�f��J�U"�B����4�]���B�6��ٓ��v��=�/��_����ޕ�.[�+��������_`�p��������^�_��A�ݢH��jдԬ���>�͞7��>�\#��U�=Ӄa�w2����g*�}��HW�%kn(Ywv@ƽ�����_8����LhN��ױb��_"c@כlJ��$�۩��o���&rs��!]�iޣv�����I�P��2��T<YK�7�~�8���2��0�'������^
O{z��.6�t>�>�Ӆ�v}m!U�;d�V��4?P�����m0&9�[ˆ�4m��t �T�����e8E?�pT���N7��ˬw9n�:�9���Q	��y٧y�Ss�J�hoX"=��Ɂ����>���w�k�v����w�+[񮻺�T�Q��vF#�H��3Oz�B^��Î�  ���<S�ާ�z�d���z�p/��|M��־�ß���F_|�x1�>���"p9 ,��C��ۃ|�M���+$�
'"�Q)�^X���j�M�^X��yY�0�d$����ÿS4�&Le�d�	֨���zp��֢2�F^�²�ɺk������� ZJ�����J͋�q�u����_5t��$Q�e�����o������S��<T��;`��~B�c�/Ł�ǟ����J���~������l���D�u��7�aU����L��Q��#���!�������\������i/cQhlm�RɄ�����B#ࠉd=ԅ��w�Ej�=ѓ�]�L;R����o���'�YQ��;m�ݸZ��
�䫗�?`{n� �K�m5�δ���H ��=]va�
�E.��^m�w9��)�!���9��;K�e�!����Ē�Պ��9���B�n��귗��oK���Y.�_�5e���+3�^/"Q���(@˚U�z��-b��1��"ף[;aW��O5g�3��'ԝu��G����/r+P�2z+�7�y}�6z�U�����{�����_!�����2[P��!��00(#dw�k��s/̗M�w=W��)��[��eJwJ�ԔS����*w��H	Ppì���j2�z�ؙ8������6�9#����E#�l��I�6]�Ŕ�j^��i�w:�Үh#&AH�z�_͢�M�Y���zo�o�3��~��-7wr����q��N6� ���4�ژ0cS�\��w���9�'�0-G�u?�`���2rV}\�col)�)s̚Ј��N!�0����X���<�`���q@ݽa8��팹sI9�0���v�=���k2�Q�L�|��F���/��
�۔��բGs�u�c�/^�M��K_Ε����c���|'�'B����B�����@S��F�&�L�IH�!�5��u��<��������<�d�ӥ�B�e���o���u�8Oo7�:!�*��VӀ��iqW���6� *��%"�lI�-����v3Gm���(�lr�Z���s�6}k{����?c=�9U��V��/�����tCѯ��2�6?*�!����	W�GP!�Dt�3�T{���P��w���N�r�7������^�K
w�W,WK�.-�9�D	�j������~k��uZ���y~�^�/p�vG�=a~�5M�I!�d �,稚I1+�WkX�_�T����N��p��	���o"ڣh ~t����~�<X������~��v�v�q�P�/m`�)���"vLBö�Bغ�_����Mq�����´L&'[����U��/�y*,^���.S���R�N�%Fh��z���@�K-8����v�#�BZh�ߔ�����_��[z)�Yz���y�R+�s�ir���SV��\�r "��^?В�k�%����u��:��Ï�@;?��-�ᚬIB�]B�ckV�i��@_���NJInJ�9�'�
><�'q'�oK"�떓�g:^�r狀��`4l'E�L���7a7V�wy�y7��'��?�O�7׺�ˬ��q��=!�����Q��?Q�{��eo@I-ƿ�N���=+OC�E���RU�1��󉊑�=Oo�R�sw~X~cb�T䏪¸�~4���Yk�ȁ� jBnv���,�-14�� �T��\1C` ��h� ��k,�4#�,�Q��n?K� ���� �&%�p�c���bZ���mf���*������Z\W��i�0ލL��������"�x��.}���I�4�Ag��L��	@9_뾇�n�z����('*N�R� W(l���A�������׽?lM
��dBwq�˃CPY!C/(�r��`��̾���y�i��D�˓���&nk��)H�����Ω�^�nC���=~�u�t�� }#�9�C	��g�9�ظ��E.H�Q���k���
W��eq��U�H,Y ZwJb�d%=��+nL���8�G[�|ljqXe���Õ��{(rf��b(5UZӽ�Md;��W�]As>�k�������¢���n^Q�U/&=�{d�JAU��}�D\�%��%2e�/<HL�(A�g���B>ʮh1�0�kHW N�J�r�˸tt�K�������0�^����g�N���K��Zs ы��U��i�e��#���zNS�=��O�A����ez����,`�*��k܈������&k���'X�97R���h�o&^;dY�$.��t�F6����0ʘ��ݳ�G�f�z<�Pٹ�n�<ͰFD|}���V�\l�N�{M	�8?���Ƅ�W���zո���ե���Q�.a�f	�xt�Gp��&��*�T�J��\�2ꖩ[r`W����,m�{���$ߏ��<��9Ws��`��eθso�~�i��"�}�m)����)�����m/s27�bc�	�vy��:ʖaC��E��ٝx�,�׬���_�\�ꁐ _�B���ա��+�Ә� ����&<�@��>~\�7;�#�N,f��.��Q鈶�9��)1�x�<����C.�~E7��a�^�!�V���}�v8�k���g�5ԍ����0��<Z�������?�`�4�Pf\��r��?�I�ދh���lF��6������F}��vl0����ܻ���Q����Ζ.�|0��1��(�gT�?�rs����t�×Y�m�`҄شcu�Ѻ��UGR,[6z�/�ؘ4�0�}H~ȯ3��G�9G\���G*�ӴV���U�$�<W�\���邑�w�( =w���xV�YD�����2��tT�F���vYʃJArW����a��u }�~OTT����"Ro$�v�k^ɜ�n�Ebn$r�z��[A�����+Nq��N�m�|��'�+HxH�����X莘�й�k:W6��-k��=DJfs�+r����$1��M��~rь�}p����{�bk��y]:����c�^��'�\@�d��D}v8����<�h
E���K�C%��o�-���YH���r՜¦���PL��/TZ��x<w�d� "����ӹ�L���{\�3G7H�*��b:˴��ςw�������|�*�@p�'� *�w���0]���v 2��]���s�6�4p!�^b��Y �H�=����3�̓j�cؙq�#�Fby��G&��͗��m��;Rqe3P2����
--朆�u02��a�ʶm �#�(���Qڐ�-*A��@��lW���/��^���zs�f�-�3�6�hP�
E��FQ��nb�W㪄uz1�����B�>sO��n�]&���A������&�P" �Zm�a�I�|��?��i�"�6��=V��p����,�$���Z���˞��%���CSG8��<W�-w /�&A=��ߟ�My�=�c�"�$`7���@���㿓�mMNW:�Y�T�
ql}�l���ŋ�X��`�&נ�E+Ѓ�Ѥ���;Bs8�Y��U�VA�p�!���zL�
h�%yT�mW	�A%�7+*nz���O7��ww�@��L�N����䤽9�q��旑�|���+��kᡄ���T?y;V���]�z_�_��{?f�Q1	 rx���Q�+?Ă�H�fI޿���=,����׸CN�N5�ʖg5�����'=�w&+-!����X8N�Z��_q�o�!=�d��wrr
rO��MX���la�=�"�kP�Bz��}���h�G�.�����,&A&H��N.i5�w��Kƥ�YN��Ų[Fݱ�46��ݹK��`�@����t" 4]�w
gY���+�Abb��kz��f�3���J�}_�8��� ��e��]��=�ć��׬��F��g��$t�_����D���?a���lc��Pn6
�� Fp�`�#�=�"�Y�_�BKt�wj��U5F.��$rVA]��Q�H�Jn>�<������b
�"_d���9��y6�.�R4No6�7�N-Qi��4�N���K#bXKle+UP���K~M����]mȜd�跗*>t�Peiy�=~�~ftU(�g�~M�s���[��x,In��9A�IE7�#Ʋ�0ߴ��{�73�l��S
������[���ׯ�^Zu ��� �ˑ�|�L������I�p0�D����~h�i�U�TS}��F[��]�Vͨ�W��Q�T�񨐄q�Y+���y�����s�l1h8	��]ً~�6l8~(�M�F�@�KF�ţ{�����k��د7�>���
���
�k��'~�`F��K�����)����0� N"D0�<8��F����eN�n��������G�*�t,#K^ǰ%j��GY�_J^z'��S�F%S�3}*���r	�S�׳�B�;�Fa�e���9H]���O�h^b�&g�f�||y����.��.VΖ�6�.�&��\!�܇�{�;�������i�^�L�$�^#�N��7m�J.}��ʻ��GA^�IG=��3�-;)�!gy����#��@�88���;W��d�;����v�����B�A$tV�""�5f���n���׃+m�e���&��i��x�h�m��؝
���&+�ok������5]�
��-a����]�tˠ�1���qB��w�ۏG�$/�H�ܮ���Ftz�Y�.�>a�mexuO�x6�r��^�z:�����r�"e�%�&�� ?Е*Y�l�W�G�N����[&��IcW��ק��ߓh�3Xf���Z����W��bQ"������ʾ�Ƨc ��=�bk	_�c�b�	�|c1�A��K�W>7�zH߰M��څ)�������������O��Y����Z�в�ɻT^�d$�t�u�v�K�@�B��s����~Z���M��t�t��\Mᮤ�.�|Y��:���cf���v���e��g�ڪq�4�m_�<N�aκ�r��g��z%-�I�8��T,Xk;.�<X~'f�6//��y�Lw���2������.
��G�w��[~�Y�ߑ��$>���|�&�|#��>}5?<�xWف���n��nwVBf��Fm����6(�����}W{|Yѫ�א�\�K���S�<��Q�A�o�^!�QUz�+'�}�]G�b���*�q�Z�ْ�4۴S�|�5��S�c��t���YS~�h��W��FpV$@Y���ݵ�ܝ�m߾�	�o�	��7D�eX�z�?O��W�gչ��={���v���^� �g\h���:R������LL���J��e 4��I�G�mC�ݺ�<��IeС�V����q�Υ7���8�F��dax�z��;�v����@S$�E,����|o����@,r������2��$�#,�!$TpW���V�u�g(����i1�[��0��3��u�"p��QcRP.O0u�JF���P����[���Yt��npЂXQ���cn~�8GR��ղ���1&��L����Q֣G��n�:��'�Z�d�ش���
Y�ѩ�����j݀�F���I�H�B���Q�1���K��:�n�ա�k\5�|'�b٢Rg=��;B������7�L/��RI���јa�~y�;����t�0��ĳ�ܯX��nl�s���D�)��x��з��>�J�7v ${�:V��-�!��9{3%���a���$��^6�d���k�=Ld���5 D%������{��o���[a�<����^䠻S c�.rC�(�l���b��C����:�F�kW��>dĔB?m�P�ܲz��Y�����L��)��R]�_�-�q��A|���'M*���`����P��嵠���/]��wê~����-��F7G@����2��e��q�Zc%��% ��#�zB~�f-��M�41��m�l�nZ�9�Y�@ǆ��8ڊT}4tŰ���o.u�f~/�Jz�iC�IQ��0����H��6Y<<:3֑<�a6�1�^���9��)	,�[k��p!i�j�U-�����qB�r; �ǆ�IУW���?�����1}1�c��~F��T��9��P��>�^�)���4�[X�M��:��������+C�!�:3��&a�*n�MN����\�9ݼ��`���xL�O�"��P�:eЎ�cו=�␣��W���Kh�djsh�Su�	�K�y �����W���c�v�ѝ�*T�z��(*����Ŀz��5�����[J浐��ƪ��&;g!��6�j~��%t�7C���۰�&C��
�y��qR��i��ߖ*��(�(�N�ġ�`�Us%�>�Ċ�Z��b��i�K�� N��Q��M�<1����1�_�R���	C�w���	R/�]��"h[T��K�]mBMg��4�dW�Ǣm�-?�q��K�L�5�ߥ�_�A��q�*�
���)��(����|��h/���1�}�@�-�r�N�1������ݸ�n���!hP���M+�u��W����t�͹ēJ����+t�o|�J0-��)���(�=(����4�ͭ�?k�L\80�/;�e�&��T\� �=���L�޷$�ǬȊr߶�c�w&�s�fiz�;���r��P��?���;�8`��+�763�(���c�Eu�{a(|顣�����Q���(�+����D�]��y릋�e'E�c�C9�%��ȱ�8z��TH�{r���~����=0����Mv60��i�iIWΉ����Ȉ���d"")Ŏ���b�����M]i�?ӵ�|�s�fJ�� 4ʝ3�7�?�_I��4�;cU�n|�`7%����.`�!�����r��.�}�E?�-1�CM���$�g��ξ�ߎ4 sz�xk��)�|�k��4�\�$ڞn������Fga&�J�/E06v�}�W�qz���Cqg1o����98B�"E���	������ �����]��ō1i߁�(Gt�D��&:���f���� �dݟ*q�p�g�2��4�l:��:�r����!ň�-Tx��vv?ƗB����RV��RRq�I�4�}ݽ}%+3��`�����;�Fŭ��=x}o�$>eh�ɾ��)���
[#Hxk�Ȱo�<��ߋ�g�V��������N
d`���c�H4@o�	$U�q�������~��z�
�0�Eh<M�c����C%ο���C6_ϬV�$��/��yutll`ٰ3�~sN_�Ɯ��r��K\�*�����9��ų�A�&3����7T�(E��`R]i�?wN|^�4�5��G6��X/��}�u3Y�!����?4���YP�E��1��gɿ�za�P������k^�c�d�[�7ݢdgB���dM�ck:M�Q��$2�Y?�N5�F���2J�V���`�<���,�f#�{��OQBݼ���g4��3�������n?'���L�U�g��$�<
��I?'�J�%nc;U��PQ����������uw�[���j�4��_JW^
� �0pR�\�4�n�C��?F-%�_�����;�x�s��!��F���n���i|����Y��3�J.�<gR���&yv�z
�9������x�z�<�Ds'(#Ym!�'� |�*/����j���n6M �'�覡U.K=D~��=SZ�Dӹ
�Bc�	+ss�8�y?�����
v��u@W��N�7��1���B��M: ��IV�f�!�����5���4�x<���+L� ���_S��V�����"Р0hr�L���zIsQ?.  �Ӻ�.� �D��-�sٿ#����M���m9���[��V�]�˷�)L蠆%��ʡ��ϑ|؛\����qޅ�K{E
�U�z��z����m�Ԙ'�<Y��G������ӟ�$�O
�z�f�����tN*��1�a�1����e����;/���Lgo\�.Eq0;���`V���2.�����=��X���N%�����M�n����Bx�z��Q����� �&%K; ���_���x�z!�R�sXK�XP���#��5a��z/�J�2-P9:�a�$�%�F�闽@Dn���$�NM���l��H�� 4�NFȋ�;��x�Nr{�u��U�鴗��r�h��ߔ�[՜_����ÏR��T�b�1u�洋����nSҨ�����Sk��1� b�}��AB�)P�����x�{��yц�������ʊ����!�^H��ApKL�NA@#����gA�d"��c����	&E��¿��=�wF�� xr�H @�kX��C�!<�(�_[$����\S �$�Bh|�C�{n�l�C�:���6aԯ�6O_���zíƠ�r#Ԭ�����PΨ RӍ�Მ;��ϩ�\��c��m�m(p���(E�'9��l�ב!U���eN����X���^�����J��n�?5U��oz(�'s��ǯ��	t�М��oPCo*��߅�R9�'u,�(RVO��ecD�W<�	)�%�s�a �����T�C~�9�`�)�k�M����3��e8F�O5��O�Ez?W�ǐ;"��J�������u[�L�e5�o8�+��w��~�u������=��bDMʿſܣ������X����|����}{vgަ�t���,(��fC��j(� hKz�Xe��
O�oR@\nM.u�Q��x��)���lbX:�?��?[G�N�_�3]y�]u��J�$�2�*aʵ�ɢR<�B腏�vE��'	:!6�ˬ���������Fmz�=��Z���� �zU���r�dn0G�^���"�����D�����p6�Iy�d�7�!���7+^�B��ļv RK��Z#ɥ�<>��H�]������.���?{�֤����ݪ��便�����ϊ�B'	zS�����_>�1'�t�I+�|c"h��y���W�B���&
�
t��J���i�����i���K�PX�����0�"��IH	�r
3<Qlj���F�̋� K���JaT����\=F!N� �����'��8�v�?�?�]�;3:aly�F�kU��k~���S��v���I�B�0�	�[��}aa>��3*�c�E����������ڽ�*�R[��5�*�'7�L�#f]sU��(!!pj��uc�l�t+��_���!����7��FJ��
�I�r�n'ezև�:��-ʿ<� :�h��&ch]R@%���&^�/�(��[�����m:��0b�,,�1tקfU�%��Ԟ���V�H{���nBߋ����⤥����[5�Pzz]���_��"�j�j�'Hb�U���*MY��m0���_�AQ���T���6�v����a挫�+����B�x�?d0�dN>ez`�u��)՛��"�jx>O�{b�%z6}}/���,+���p'?~��z>�҂�)<Fz��!pz=axu��='�T�EyeZ3Tщ�j
 �G�P(�}���Aɟ)Wi���Nޟ�C�cRw���%	�6ճ~�Z3Z�0H΋1תe+�]�d�G�m�UU�j�5j���^E�-J�����ڱ%%�R��{#A��Pb����f�u���w)t��ϟ;y!���&dQ�(�/m�>����&��,Hc�yя�O�L{���D�p�*��.��h����� �s\y,�W�� ���~�}��;�1�F����w�/�}*o�Cq*�LM��6u�	�U׎���B�E�
��\��n^����ueP��Eyk��)��6�Y ��&���~��
�t�r�fk�x�ظ�<�6O �����ص��3����}e_k�nz� !�q[��pu�9ܔ^=�<۷�v)�ݙ@U���͗�D���ShYs���M�������tI~��A������1��R�Kb�!5}�i
 1q��޳ޒ9����=�Y�b �JmCAˋ�j'l����|���?�DZ�p<Sˋ�f���{�zŲ\8~{�Z���M_��z(vi������4z\5X��9�Ll�v�꬇�$�� '��D�ď�!���+u	w�8Y&�.g��cb���`���!��^c2�$$�Q!7?�1ʦRl�����n m�WU��'�S�:��������-}�c���Eý���2]>jV^�~���t�ъ�wx�W�����D+މ���α�h�h �{H��UL�!�%e-�����caIqx9�]=Ժ�i�J���������sݽ�52<4�}� � Dt]
Hˬ���?+!g`.T�G,^��di(�J]jyru�Y��@jv5�֣bې��m��$+�6moZ6�ڨ~� ���f�`����A{`�k.���
�����N��|c�g��'xm�s���Uں򍁮���q��5���=����K~��)?,<����@����e��`ه������РQ���6�f5�寚��˧�6�n�"X��Eo��f��C|��I�b���|�T!Z!�V�9�'�w?���F	 �`^��<����q-�]��Eo��{a���W��w!���'�������q��J���.Ҷ�/����M�WJg�3濤(НnƖR�*'g8ҿ�p~~�A��:��%`'S�h�c``aq�p��<dy`�&��%��R�-`t�A���DhǱ=�Q��
�����3��Gw�Hv��i�(nא�Ժ�9�M�A�0;��8?�fzO<y*L���S��~�F�ϲ�`�n[h��,��!_u���r�:�*3h0�g�q�e�����.��(�^���)���^�$;�kR�{O��k#��Y'��A᫹x�O�P�h�2gӹ9�`v�G�8�9�he����<�-���tHs�࣒v#�HQ���8�@+,�D=^�vQf�O�m���|S������s�(��O%Wo���S|�TyƵ���Mo��:y���ھ�3�R�`u�  ������:�'��6{��h�N���`�M~�[=��P��qA�e��..��щ}��`Wz)�m�{գ�v��E�U�ǽ��u��\�/�d��2�����ʹy[Y���Bn�fN)+�8tp��k/
e�Ghm��7|*o�ڈwǻ�b�d?��S:�����ť0j$�Դ�++���O��tB��f����p�Re���[9��~��cNE����m�)j�_�r��wUU����h�*s���O��ѿb���,13b�gƻ��5bU�d��I����?��c�E]����K+z�QB�5�O����e⮠���6&���6���͓E�m;���p{V�ޜ�Mh'�c�٠����;��j3A���@f��yz��T�%�c��Ov�)�;t��t%���9�) v����M�ju%��F�rh��	Q4��:�;�f}eԏO��\M��50�nX��c±F�������i9�H_`�a�5�6�0߱�t����ݾ/m��N��Z���g��l��6Ѫ��{�b��E'���]�OM,����=� �����Q�>'��ш����<{*5������Ƨ�9jj�,/+���e���_�d���-!9Dj=#%�дSmæ�t�r���2���"i� iL:LL$���u���7=��O�~y��z!`�4���r��.�����rJ��ES-�����ɳXFZv��uk��"�A�� �C�BL 
7<99}$��Ώ��׶0+&׌��ȷ�D���I¦4w�e�l8�z�'�f�	�چs[񸳑�H��{Je�1�M�8�9]ʘ���9_e�d��{{g~)k�����R�)�j��iF�N�����e�c�^���c�mz��x���ut�ƾ�I�v��-Z̥�[�o�#.��D�&��E�G��3�/40p���F�8�.���F�~!��ӯ��K3�o������E�\���f\b�5EewgW�G9]��8����;72�U�z����k��)3�?�������)����n������W�~So�>�^j�y�r8ߩ�1PƤ���vTl7��{��hA����f�y�(x�m:w\�?�7��G%$`3��ʯFx��C��O�u��a~U�L��:�t�O`���.�m2*9r*�}P��9�a��i_�6�>Y��ȷ�*3�߃��!�O�ʼ�>�wQ��N��q��euTo���L�\������Hm��K�࿄�����P���j�e����ͺ��;a��##�&HG��ۜΙ�6�V��]i��Jཟ�j�	�ooj�s�cAh�\]�3���;��;�(�:4D�Ngt��s�"b�`�.��$3(��v�ac����~��
�}ɋ@���r�O����)��qk�kk�Ӄz�.��I\��suz����Ao�)�'��ǾH����t���`� ���fZ5?X�?7�_��=#R�__�oG�c;�k��o�t���@��t��凓���o��\�Ic���Z\;k-�$��
q����ʭ5�/]�n�~���w4���1J+R�DP`^�t��8���d�B�|���,�Ϻ�`s�Ųv�׭E���q~��$�( H�M�plj�"�L�M�
�0� =31��<��������KNڇN(8%�*h�5*�[㝿�5#'	�-��Z�N*֍�&�k!�M拺[��)�spη{� r3='�a v��^���'ct�Z1�6��I�M��*���"�Z��9�$Ų��-Yr�N@UU��쿟�{����|^��@R���D�\'¤ݨ�����Yc�AH���,�!�����;�t E����H��	]o�tޏv��w���vq@�-��M����f��	�f�X6z��S�Tb�s}6�������C*���ٞ�ȗ��#�L���E[�>�2�Y#L/s &���^�ϡ�l2gg�gwL���,\eG��R��j�M��#�XI�7�]ܠ�c0򿺴�,��K�,6��ox��"��Ÿ��p��NDq2+ᡰf#pǭ��R���IY>�>7��'+,o`��ގ��+�f} C���]�H_����q����5�Ǟ�#�B\���)l_��f�$�ig8���t��p��ɐS�tZN)d�xw�J������3i��)�W��H�v�}/�_�(	P�L2ͣ��GMla1�O T���o���lB/�%q4BuA��2%ɣ�]k�ʴ@6��%��)UJ��ۋ#���r}=�O��l/��"���96�X
_zD����0P^A����vi;Nֳ���+� @�/�W�6��GDl�C�؇�;10�ϝ�y�)���͈�/�05�ʬ׌[c>����'K=[���E�VXT����� yUUՂ���j���8. ��S�)�:#���j>�a_�k+�i�kC�0��|3�@���`��L���>�!���Y؛��C%��V�;�5;GKf

;��Z[��R�����ڣ�EGw6� �#ctd8UM����K��@�w`�0vq�Ou������2}�؀�)xK�A!h�J/t0SN��u�^<���\#�G�	�(@�M�}�Bj�﹗���h�Hb`��Fu�����/G����7�,��mSh�k�O���/��<�&|w��srnz9v!n\�X���sq�:��1`0v�+���\�U�X���d.�p3�M~B+������C6X8�S�y��V q|��u챯�=@�j6���9����eB��.�@5��d�e�}Xβ�|F��ʸ�P+M�.���ϟ�m��Jny�J��L��M7��ED�0/���oMNL���
^�F�C"j��ǚ��ow*��(T�F��Ýy-I�Z�&Elw��d��J�ꪫ6�>�V��>��wt�f�F��QͿ�<v��ck�^���".n$�U�`�����{_݅IR�
E�l����W!����Id/+�S�J��*�",��y�,X�q��X��#�wRu�.^I��%�8�.�j�e��S)6n|���#&`����#�����k�oaW�� ȟ�2�l��3��R�r���a���J����W��N澭�aO���+��c�R�Kb1����H�q��C�߶�_�@�rI�ɩ���9V���(��7O�x]K�=TL�YX��~�;.vD.N�P;�~�S�X��?�Ii�Ek�mj�B��o7���$	x����=2A�k�M^�3�d��D{�_��^Um6��Qm�C���87�:�mH�ʗ�a�(Z�K,yɣx�@g}����Nws��p>@��F�o�
��S���5N�&��5ԔՑ����/�����h��h�[��.�H���J�щ�Qf䞈�S�ָ����Z��Ғ�统��fQ�[[9���((y,��I$�>��g���oE'f���z�p��o3u���߯N�ɥY �3�&`- ��?c�	]����vv�'4'��?�}�	���g��jj��i+��\�1��dHH�r������p9���2by�B�1�}zH%����(+w�Iw�o8�}C*m�I�Wb���@���Q�y�7AX!�q��E��c�T,�:?lr�!G|潸�VV�������2Zy����nq/�!�qԩ������N�������na���T�<��	 FJ��������v�q��_�F�;�-��S��)�`���w�D`a�! ��w�����T����/�GL���[ف����A�
�����O"�� �$��:�52���
P�l1����$���)Y�p�P>Ars*�lܿ�q�ݓ �x�T�,8o'9�B'�&��O�iH��cI�b�;��9�W"V4�><,��B�v�N�cwT<uZ		�)wU��l���|'����dL��QiDR$�4��=�koS�����(�l?-��u�bۖ�P������F�,�,��&��j��?Y@3�`**k��e6�hl>�r���?U�a|Zu��#8X2v����"Q�r�3���N��\�ˇK�./�YF�!9��켚��ˬl�BW!��v9�u{�o;ͨ�e�eR�O`C���p[N#�R��@�7��]�Q����*5�^�VHE�+M����7�냂*f�rsn�!� $#���V������[�%v_~��_�/4*��ԙ^qN�2c��L&��ANv�M��TG�J4��3�G��5Q �u����vp۬o�Y�W�i+��/�f��5��G�ꟊ�FYUW<^]������1ʇI��X��]2�X<��I���;��U�2�]=�\�E+9l��R��Q�X�/�;kDf-�8�bH
�p���$O��\#�����!�.�ZI뷟5J�� ���F�Id��2&[��SZ-dx7�J���l]�[Z�bR����5u	' A[�����5X��Z#���+�� ��cԌ�|�:��]���R9��nKB�}���L6�D3_����t��P���PY	���3��{��M���������p"�#�pΑ�=ϸs�w��{<���>��x���u�w�d�������K�_�#���j�X�B�(�����S{:�h��'C�À�P�]y��*���2��M�3�|����_`9�]��|�n�n-R�Lg_Z��ly���*�^����+Z���}�*=+CF���B��$|�E������)�Dཱུ�z/���t1�����=2�o� �>��R���~����Y�{��
��-֠t�_�+GT�7��c��E�xnQ�����'���2����4<s��j�Vj6��w7qt�� `Bx���C�}Q����D6�Uz'G�X��âu�-Y�8M�MZ�?��7��3�]�ba+�/��_��K�kdh%U��{&��&�x���Y}�J�.e�XKeg?c*{Ŏ�� �&���7�>�A��I�R}���W�Y0����SӸ�{����[f`m����q����mCA��];ԋ��f\"E����v��,�`6���'�2$��b�/�#.Х٣���%�A;<�@T�j��" ?�������� @���ʏ�C9�1�W�i����6v�ͭ�>���D��azZW�"躻���nb��>�7��pK~��˽�#g�=�v������:9�Y�X¡5�w�[���)1�@G�=` 3d�(�T|G@m��`��r�Dl2pp�<Og�{�8t���V�>�W�_R��ϰ����3"�0��C��C�yt'w��*�)P��[D�� ��??��q��|�uW9t��jQ��~��4���|�<Yc/¶�ZS�n�h�Ů�*/��õ�}����ty�xP��Zf�|�8v��|h�����Xr�CmH���p�����$����(ɱ�%t�S�4.�c��$y�� zZ�|Mӱ37/~����
a�`}X|���JTD�xN��2�0=�I�0���u�W	鮊���~=�	+Z�B��Qh��$ο��˂�Χܫ��Y�O:���mjytvkc,�5��~���-��;�զ��RUf{Nz.�F&�]J���i=�if��<}ZRBIO`(A�feY0���}S{V�E�(AQ�	�E�+�D����A-=U�5/^;5�r<悽4��O�3wi�$(�>x��u��N�����ƾ\�V��� [���*�!�d�lϦp*'E���������)'�%���ſ�N�@V�� fEؤز���K�ۃ~�u{�?/�e%(��gѫ|�L�Հ���J�G�t�+�q�Ba6����������,�ϸb�-7��2l��,��\���`��N�� C"�'�M ��N�h�鴵uw���!��U��:���3� �~$��W��Pͫ�t����Hx�mp�ޭ20W���-h��ca����c��X�Ux�d�+ڗ3�]�4l�'jr�]ЧI��������7�7h2X��[��ک�TM5�У8\��!�
�3`�0����=�@җ����Iw�y��q|��8���b����2��%3i�S���c������H>�G>�ЄUE㝝Z�q�����~�%4��Ф	�e�l�k�](��>�2J���+�0<�a�<�G��A���g{�X�`i�E��.8��.i��V�'_�b�-�ɫAE������w�x�&�q2/�M����p���ަ����0�������N�1�i�IZ��:A���
`��g��\'#���� t%*.6�
�^�ￂ���}]̴7���O������zM�)�M�{ܩ�ּ�w[T���ә`(�ү6��G�?��Ye��5������I��.�ɨO���M2�*���2Vj������`#&'��ܣj�Fqu�w�Y��JǤ��޼���l�/�; Äi�P�G�cA9�ȑ��/�wR^���|k{���(�}�Y����}��G�
��nF�M���V���o���9|��\����]	핣�68���0����"�<�5g��	ؠ��'�S�l۴���9	��졈�hX3�2h�7�B�O�g������������?vO�o'���qhE*������{uΞ�I�AkB�u+�FB�xٜ`��z��p�F{8�C��m��\�(+���&9����]��B_,�xSN�P�t�#���w�.����݁X^���G���4�YPsoC 7������Li�=+�XV(��D��~V����q�1�u�I|�)=ٞ%��|:�m��EЁ�ix�*DR���#J���v]�]��%o���t;���[>�u�e�tx�;.��>�@�������Dd��>���WI{�	+޶��Љ]-%B���{�*dXĖ���d�.ۥkh��o/�u}�n�w&6��w�y#�|6�������]�����o�~�m��*��'*�6)����v��9�*W�-)ÃX��ق��{�A��־�/�З���[�l_��&(���n��(\��O+$ﰪ2蔝�*"s̓��H;��ow�!G�����9*x�����_��G�IO;� �����ݭRE��\q���xg�T����/.��D���l���*A��-��3�^�������%�.x�eV��Ʊ�d�w��[[+a�������#��R��?�+�z��O���!F��ݩ��4G~��r^��%T�	t��`�줮`�������:[5L[5�7E).�}G��w>����4|��۞y1gl���e^g�"(�1�� �f��o�� �Ɠ�
��ea'{�����Y�'.՜[c��C?������
�\����y��>N��E38A�kw���zY�D�z��?�)������ڌ�s�:����3ώ��/�黻M�����Sݻ��eL[c~��X4�>^�.���eK���j�o���*
�1���>Pv)<_JR�D�z�y���+a��7��������qq11ƙ��g/�ƍ�"�
�Pa9���k��3>6� ��g�wo��������v$^���.�׃���YW��adaט�<�"�zo�� ���M���8&N�fi��0rI�ƺ�(>�TxϤ�NO����}�pK-�ޏ�������I��Ĝ0[�@��jcz��˧�o�q�Ww(CL7�#c1���s
C���o�+�%�M��Z.�<�`�/����|��׈�����M��o��h�.w�#���m�b:;7�9z)�(غ`~�l䭌ȓ>�'�`��^���w-(g��K�&� ڲ�	u����@�W���iH }�0]��I�0�u���	)BЗO-���|n�����@@�nC����y���Tp�|A|
V����w�zy����k��Z���ozD2������K�>J۳Փ]�7�wHr[9I��nچ}���rUo�ֆ�����V`��2�[���?��z�����^��*��?�,�q��m�����a$�MJ8}�m%\c��uy|o��sĻ��.���l�>�Vͩ�*�?\��ܔ������&T�Ð���`��~��S�������;G���O�ji�](�ܨ�K���&�/�%R�ё[d�S3?)UNUFf�+�ũ��	[\�.��O�a�c`�J+��v\��Y�R���ļO顺Y*j�5��?����Gi��E"��=�E&����h� ���a�7��N�?sڣ}��H������4��/}�k�|�v	�n��T��w5�7�G^s��D)1T�|>��誧�f��KmuW=t�O����şf�%��|bO���ɡ&�̡dp �Q9j�����p�b����
X�Xb�7Waf��̦u���9��S܎>\��ɟ����恼p�"�<FrF3QL�S}`�xa�un��g���J�����)��^���������?o��e_ؾ��~�tl�;D/�k(�c<�QVe�i,�z�Z��'�����]a%}�~�TƏ����&�<����_ڜ/��{b��A���.��ō5[:����+��!����?��� Uq��'�
C��6��{�w)G���0�(4�G(|a��.�\ߑq���Ԑ\�w��AJ�>�"`�7p}�VffU?5v�'���������=*k�?%�f˭�D��<�vA|	������몡E.�����t?x�]��`?C�`���5٩z������ܯ�'��ϰ~���K�N���@AO��N�kaa�P
�f!5:��d�{������.��Z7�����w'����=��l�U�^���"=������G��iMi ��gr���蘑����~����R 4s��g4��:�5n({�E�5J�:���ȫ+!#���^k?Ѵ�p�)����W��:�*Z�G�ܴm���s�%(tn ��I�Y�K��Lt�Q>�k��-*,n~1*���`6ޯ�5_[���cpȤo� f.��ͩNKt��
��0�u��,Nmg)��թJkcO����=��9�zSb[�Ta�����G��yăz���2:��&s���g����.:�fY$w��;��]����x����6o�C͸�=é�p��مcfˠ���"a^�l����N��%p��=��e������(��[�n��`�߫���	*g�7�8��(���$��˦�E���h�����h�n/������/{�`v�6�,0a>h}h���Z�;�������ƚf5X��ib��>P��t�Wj_X(��0�+�d8��W��x���2�,�K�.�g������(���d���2��k^^��p _�-���z��8�w�G�?���ȍ�c���@��S
��aWk�y1G���k��p����U����Z��:�D�=���dd~H�>b���YO����I�&n}��E��K��ո�y�ݥj�=�ю�<ߝ��wC����Y��p���}������t}X�i�ӕ�ޞ�:� p��;��Z\q����oѠ�����=ݷ�ǽؗ��q{+RS��5ٿ�59cC�]��?�g���JLlCR���g�'�	32�v�����뒆���FBş��?wT��u� T�r���e%�:]ދ�f`��M�^U�P#��r�%4�}����	�"{t+����V�n�����^���+�X}ǽ4��ƛ�I�X)�P�;�Z�D��������ǻC<"	��N4�H��x$t���RrR���Ѳ:���KK@'�/�Z������A6ENQ�*/鰍篞�;��=�q��x�1��ϐ��_S.��j6���h�N^6��Ңp>�m��4�K��>�.$���d�imn��x.bM�;Ͷ򘞧��4f�lv�=�&������D�I���\��I棰���-���gG��R� A�mL��)��W���;:�YÛEA��T��g�)/��%�xy�{�M[|��/�;�4���1p�#mB9x�t�߸zMr1߶yǃgM5�J �<�H_^+yU�a�\ă�j:1$f��w`�2����� j*�W�\D'Z�O��?�~\��Mׅ�^T�S��Md��Ip�d��Y��iu����s�J*r�E�4iJ*ܛvf���Y5n} K;�Z��Fz�b�dM�i��-`��.�D���rE�p6I�[ I�����>��\F������}k� L��(��#6L�?y7�m�Ǽ�h�hw�����mY"���d�������P��k��Ag	�!p��ySh��b�Xp�N}�?���}�+ߤ�����BV���I1�%�\�V��[m�mh���Zh�{C����Ѯ�A�.�����u�s>�ֵ;�{�+�k�c7R�Iǣ�Y��5�ۘEIl���}=[ԬZ��+���Ҿ�F�.@bB/0(��h�2*|���wv��/�軭W��1�=g�Gq8g��	m�ޙs}�)���.��ȼ��W	�u���������x�6q�x��]3�<�s�)E���ѯ�,��9���GKc�Rz�����OG���?*�M���+�A#:$t0�Ц��8���`��T����FhIgm���] E���*���b���A�UF	h��'o�����*%�v?��<b��ǩ��;�Yb�V���h���_��e�+����������QI]����7A�J���fJ`���Y�w=;:a��1V9��:�G��*>��&��m�%7_�;}�oe�W�	��𠥛)4
)$��Ф��4��oP���ëd�9����}��6�︾�~ %��Z��m}�,f�$�Ʀp��e#����j�$��G����0������I�����ί8�R�GaA4�� �'��dx�ڠE�v��pa��%f�Ywt�T�ڀ����_:������=�?혐�(���6���������TGr���ka��)�d���\Ϣ�j����4�ʭ�;X��C!]�6k���+��<:�&jrN!�[S���_L�

��p>?��E�&��d��[�`�Ub���H�+���p4�y�Uc��~/�����- N��\x��f��Pl�U��+SY�V��.�)0��kp�8��ۄhTI)��ʒ��~�vi�}MJ_N^(�;e�� ����{{"�?��[�#9�6f��hut>�]��x�x��r��|JR�1/1B0"(A�U�C����;p!}EK[ze�X�8	ߚ�N�ٞ�S��J�lo�[��&���J#o�\U�hh�.M��,a���*)�4�;5�g�E���D���H�:����9hU���Ħ�{��s�]$�ϼ�q,)�����ſ��M���\*�_�@@��UDM�x���E]�V���<K��qRn��,\�߯�l{��V7�
�t�Ē{\����
�v����(��c�t0)r��7UI}x�?�w���Er�r�+Ӷ�|�@�z�Bs8���U�v񌞚؋'k�8>?[�hJ�#v����`5��Q��]��lj���_9�M��`��a� AG��$P��m�X�k���zZ�\C�#�!Z#��N��uH`�����qLf��jdWhd^��u�e�2�=F��ǫ?
��������r���⳪�,-4w翐���El3P�6�~�5X|�	��~���մ����.7�R��͏��\#�{䈀z,X����s��eS��y�����B�b��h��BK�|;U�N��O׵K�j����?:�z���Ĝ�Ą����3��V5��m�:��3BY]��<6<���q��Rxi=<�Zu���D}ﰛ�"��{�=��*VG��3]NcK�İh�܀R�el?V	\2.|ߵv��"���������!��
���:�K%�g�����}��ɗ��q����\�����*k			0ә˿��_��ߢ�u ��KƗtJ"h��_x+~�v��U���S�.�6�<�v���v|Y/�1_o�A2g����-N���HH˚E��p}�82�N���ޝi�A����t��>�9�o�#x�N�7"�,g�;$�\<��X���<c������]�6���s��}Y�_W'������0�!M�N�ND�moOn��&���I-���O�ߡQ���n�U솲�H	����Oq�[*�8��>�H�N�6���?�k��c�z��؀ix�߾�%�A�'Z�>N��&N�S��>���.G��|�U�,8^ǪJ���\g�65 )�d8���u'�G��를��q��>���0���,����b@Q
4�	Z4���HH�ׅ��(7�����p98d�s�Wk9�۶�^�>�cx�3R����FX�e��0�¬�4�17G�}��`��P�(����bЉF�0���=���B�:gJ-	~���j;U_x�[����{�1��u��/������4���&�N����P�c9�t��w��r,_���L��O����+/�Չ�'�l��yJ���M-p$F����E� J;L��#�B<���yu?�U�?�����0�\l.���,0dI?���6).}ߺ��3�1���ڇ�GNW6�OD����C(���x�$V�Y�<���P�|sԕQ��?r��k9/��j����E��N����t��G�FVW�-��z����i-"c����b��Z�����6Ks�ۧ�������TY�9�;a�G��oES�v�̈́s�惮�d�A��FZ���ӭ�D�Y�5��ce��dc��?|��h���\|�z$%AO���+U���ѡM3rVz��������l�Fuvܩ]�;�!6�ָ��X����G9IޥA�F��:���l:@L����x��xs$j8YL��(Y2%raǿ��;�y'�g�����l=����󇁺WwxN6��9���<Eo�8�R���A�"���>���x8��/��z	���O��ש�N��Kڌu�S�����\bf�s[x�5�Yt��\�윟�2f�r��R�&��SE��&v�P�]8%���H�\�����}�d|��rߧ���H����-�|C�M���G)#�߫?m��2��E��ZCbK���*��^2孭�2K��%)եk��k	BWۦ�_t���e����a*w&���C�O�Ţ?�!_���ܱ�=��?(�ݲoʦq��@��J�=��2��uԟʋv=�@-y�i�Te�6�|L��$�mmu��U�!����6�{9	8!��z�2׭������w��>��#z"�� $�4J��Zn.��f7�"�vY���91m�ds��i�_8#}��Oc�Dg*�KPo�e�H��c�F��O�:9y��~�^���%X���;��BT���W����_|k��*J�j�l�g�G
���M�G�H�������pE�grmI�#�w��p�{�y^���yyٽS�J�� ����4�y��wf���~�ߙM��m�-��z/͂y��7o
��+��i[�z���|�݅��1=��O�5�MB��tO%q��ǒ���A+�@x��l�E@޸k�6�����8�g$}ٚ�f�I��ː���~"�'Y�I�YN���=v�@��Iw$�g�j�!����=hI�lo�VPaa���2؇�
��˛A,U�n���^�mN���ڛ2�2�c=�}J�it��;Y�%�34z<'	�09��Ly���^c�c���N�֔�J��0�T��Pg����]�W�6#��g��T��������kA."�������
��N�Cy��-���_b2�k�˾u>e�Y:YzOԭ�9���i�$��f����"^��k5IqQ]��X�b�]���U폩�￯V᱄r��n�e7�x(0�",q�I�~D+���t���
��2,��_޶x1
h��"s�˗�IL�#v"�]�/���>�~ۅ�HD�T������%�*�=��{�ft �3���&WP0z6�hl���1�$�o!)��Y>V,vo�x���˨��Q�xdRk��P���q��sE�wC��Q�TWXx��\U�i��S���A:�`;<N���15��k�N�
�8�2/����+yK5��+D�.A�55[%5�$%�!A�Ln�I���<jƑ&v�*��a޼��
~��,��Y��g�[<�!�3t1�E@=���5�}�_�@��Yf���X��痭����*�����nB,Q�G���0_ɣ�����w>���ѬWI�	=C\p�ZM�|'�`},^?�+j6�d%�_�5�c������S���*�7���zmm����:w=�ZO��O�?�{;���ܣ�=B)(�F���e�^,�9�#��ʅ�
t�����OMcK9݁T�]~ܾ�3R�4�
]{�����e��T�=�"�p,�� $�t�Wz�?�K�]�[S��VR2Ȭ�9Y���P�����e�S�H�o��.vO4���e#7+QZ�YS9%HAmw�*:��F^��x��HJe��^�t"܌�NJu��25X��<�w�K��'��j{M��M1q��I'!/��I/x����y�b��*�-�G�53/��U��s;�L�.��_p�\�7#�׃��ot���?د�:�� Mt��ׇ�io{��@���0���{q2X�3g8X2G�3�	}7� ?w����R	�'� g��$w�׸Z����wV�D�z�gϺ�-/�_ױ���KV��ؘ�mJ
}�mm:�+5J�|´�v�P=���U������Di�L�tiC�Z����u�E`�39��l�sM�Q��[&V̪$�����.Ɲ��._n���O���s6�@C���L�z���ȅGwE�&��҇?�{?�E�_A���'nr���>�@.���l���1�r�A�f��f��E��q��W^�O��3�q�Z��i��^�u>����2[+#/��xnC=2Mz�����0���������5�၄ěU!��*Q_|v��'ʤ�و�o
�xW�X�b��Ƙ�{)�υ�;�>#ڥ��U�>���6�82p^�u����9�� �&(o�9���z_��D���9#!7�]����d��$2�߲Z���Q��|بLug������4�r�Uz���M糳�kt��� �t}x�gR�P^n�X���;L�@�c���Fڑ�O�����6����a�����t�jL��K��*�(|%Pw�����%<��U=��|��S[��L�_|��?L�%8�J;+/�����! �����*d՝�o}�t=�3�e��5|5�x�yS�׶�x1����������tu����Z��ۗ+��}��ج�W�Fu��<9:�7��}��0�x/�T^��8w�)f ��t*�ٝ�v�����?��W��6��l}v�f�].��͸�ٯ�ỳ�����-��߾O/�-��v���3P�Q=� o=�
8�-;�6�b�OP���[l�!���d�N���ǲ6eɤ��]����r�iE�1J@[C����	��t��G1����ݹdl�(4:TA 17��?��`�|�A��m�
�F0��wC,Aҹ��xӧ�EѨ�X��C�0�}'��}�	�c4�Lã�ǆ��q�����%��a���GE";�����G���r�)#ؤϷQ��K����ف{�A���VK���z��7 ���l�L3�a,[!��tV��賣(�uy�-��i?���r/���^����u�2�]HA_��q�,w'�@��앤72T��MWN!24]~L���2;�?FD�HfFf??|t!�]r��,�J߼}�&��nzp3�Z!��#Oy�OO�C��-%�ٟ @Ǜy��'S��՞	�
L��	r���oo�<.C��.���9���u�@��%=��{#�JA%��~��TP�6�:0P�b�����1���7.���$6�+����U�����^�o��?N�0�̎s���U�G�Qxh��G��9V��e���!�'�Ex�*��F���	��i"p��u�T�k�[2������F"[���;�#��:%7���7bs$"s�"��Sa^2Znp^�C$���󰛯-�\<�7�à��������YϕԆ����l��6>ߥJ�	89u��/U������;��[�̚�ڃ�\)��Kj/�sa�q"aa6�@�^k��4��\�n�q�e�
��d�<B����촯�Z��-���nY!f_e��%3V;�]�L\Q}�g����Y?bq�:�oŴ�,]A�/�Z��~c�y{��5���P*tM\�Ȃ��6��@����GLz��j�x3}�BԵ�v���N-P�v�s"���Vt�~��Zǩ�x�p��n��ƕa@�#5�H���ud����Љ^��i���|�r�^Pea~U��0�������}�O�7Đ��&��d�u}!u~Ѳ_"�?�`��Hf��9D�/�3<���r�tH	����*��T��}��������
�R�!�099�{��Vx���ٔE����,�]}��;5w�C��߽Y4߹�����y�;s	zZQ�i4ιN
Τ$S��i�2DȔ�}C;�l�+*CLQr%*m2�)��>4���'�L�"�z�,2�����T>�]~��F�f˯��]�1K \�%�T?s�d��6��&��`*w�l��2P���q\��fN�P�"��J�E�3�P3h���nҫn?X
i��t`��*��k| �\!��2|��|�8S4k*t��W ����!���E�*�u���;�ޛW��=h��W]�Z�P���Q"ǯUދ�H�6(#�o�N�.��y�-�C�O����\�C�߾�b��0^,����-l��;N+`�t�ɃL^�uS^�s*�����z�
a����o�KLgp$�e��pj�(�ҞQ@jM:	\U�=z��_>�ŘfL�%,¸YzZ+��i�tt xǀ� �����)D}�
�;�A��l�M�x(ω��Жmrv���K�~'_�%-M�H���X�_�NQw�+�Q�
����l&<K{�u��Q�Ժ�.��>��Xk�j
������0�\Ӗ��Èo�m65��"���Y����eͳ�X����N_��W���ʰ�7�#j�g�X>Vc����^�]��}P	��U���a]w3n����|�b��#�P���x�?��Q�����%��\�Ay7�8xfy"���W��e�}�3⬜*�G�mm[eSo��t�R%����X}l{�s��)������?r�.r��F5�ps�W&����:�z}�k�බ�[�W�"��%*��I�g���������kk���Dn�`��eʾg`̐wF����7�$`_,���V�����H���~��AWoQű��pV"�x2� E==��{�`�_͑n< �B�:�_��B�kj����o�*%p�3N��cNW��!�$�?�a9.H�v����H0/x�\Ig8u>�#������2F��> ���y�H~�I)�h���J5�Us2^{��v[2�{s�7k��'�
F�l7[z9�X���@�ܰt���Ga��E��C�x�v���$	oO�H]���J�רt z��(�,�O��K�)6n��j��m%�Sc^jg��}���eĥƺww�hC�'_�C�0�zJ �7��!"%ƕ�l+�l8U�����v�K�G/��&���FN�$t��g���0��<��2���0�p���Y�����o|���0,�<��cl�Z��;�<Sr~l�A�,W?��õ�Ϣ�d᫳�3>�sKo�܇nz @�k{�gvpf5�[c�kݰ&���vo]зi���8��k[�Q[ۤ"�~�Ȍ!�L�:.�w7�U�������/�%k�������_]�xmBlZ�8���P|������x	j�M�Z�-mѾ����ݩ̾_hK�yo{�>a$�ߊ�8_���*�iH�܆�R�i]��պ������k�%Zt��*ºt5I���nxd����N�!�����X�^uf�E1i�N��t9쫁�Y�3���jﾟڇ��R�v����H$c����ɯ*Co���x3I_����9����������^�!�ս�=#��H�B?�6QF#���G���i?��@�lCD�<���n�j���dɌ�<i^~d�9^c>���FL��H��ồ�O%5����6�Y�A�5H ۋ{SA:��';��/�l�����\}y���;]�l�1�7��Q���������&Oe�&C���������6�"@�盛i1o�o�@�&�Ȧׯ�h=����X{9�������)-�`o[h��j�]�1�^ۈ�6ml��<y���r�
��USG`E��0�E4tE��Ǐ�s���2�l�V�_��G�m��u�/�@Y��KS#t/�I���'�8��$��3�C���@�Fi������bS*��u��GKzaw⏟��;�����R!�y�y�dy�]�|{�D;Ň:\JA"�U1B���~�5�����ą�zs�5�)� ��әk�"t&��U�f���&��g�	]���VJ��O���'��|е���qF���ҕ����`Rex�@���W͏����R����� �%�iL�/��sL��)��`(�����긴���׽�QX����\�@�#��ǡ����K����Q�s���o`v# �㭠Cf���N�	����׮[�zܓ��c9x2���a�V�ƍ��r)ۛ����s~4)���갅E+�Wǆ�,ڡ�V��ⷯgƹ��?�SeE1&.z�;ݮl��OL,��J�o�]///�6H=���`�])�+v�m6ǿ��xyg��wG%��R1oO7j���X]�y�܏yUR�\W��ϼc��̼^.S�l��<Ϊ����ȧ3�JG�F�����5�l��}�D�H��]A�����i(�$`d�s�`e3��t}Cek+E�X㳞2���%���b�Kl��y�tv����״�&�x���!J�~-;�Tzw�[TL� .�]�}�if�A���_N�1`��Tr�T���S�yL�c�-�.�L��ᮉ&����<�ssys�����렑-\���Y{,,ݣY�l��h��TiFn�e��X|�d���ުj$��P~$��ɿ�p��/~���Ǖ����i�,[n.8?��BT���7cQ�����	g�5���%�q�)5�k��/b5$�"���{�B uږP���7)����	��Sh��G$�vT2�'R�꣆�l�;9M��Y`ob�z�ˊ��Nw9������h"ո�{w��XQ���d*��0_}34r`�*#P[,��ɫ�X�׷��
@����'��Jg!A�0J�4K�G��\��s�v���7���~����S0g�i������O��LE�P�M��`h��@��J������,�0� ������O��/�ixޔ6o���8T&��M�×=�G������l��������5�N���]�h�'�.���1���ɮ����p�*����,Oγ��.�fba���G��[1hlmM�8�C�a��PK��L\��[��2��#?�=��M�a�Av�}/|���������e�M灠`��eq�N�Bn������+����bgEz��÷ƀ�YӍf5fAĶrYk'�&9�M�~o��O_?�:p*1N�gg%7b����!��d�8�!,4U��<�i����	_�'���]�;�D��<(��k:rԼ�{�v�>�E����c�y!Y
Ģ���(.�T���+/����[Bm�s���>+Xi��-R)����;=�����o5Js�i�Oj�G����i��k����e�n�ҹl/��"`����8��U'Ř?O�P~S�?nsN��	��O65��ȝ65�V�F���7I�f�:촀� ��	�a Փe��5C ;%�	7?N:���:s 0�V�W��g�h�
#��?qU�K���rv�e6yX"��B}�W52��я ÓW�T`�s��Ի�?t'^P_�·�|{�ᙃ��Z�sý����lyy�͕G�F��j��]|Ư�rK�}�[��������Dܟs�E��~��,)��C�z���z��S~����(|7�w�dcԐ�
p�xY/���3���?6����Gø�W��.Y���Ifa����GtK���6}X�̸�S=�qWsc�ΔfI�x2}�w4��Cӏ�T�;�'�+��F��}=����gK5Y^��Q�V9�rK�.��ю<*~�y���A�!�R��HysD���c�G�]�����Y(/NimS���A�⤴�Tpf��H���";����4�$�*~��dQ	�����zU�?�SM�����wB;RsĦ�X �̯q�-�+�[�/{�3�ߘk�q��JՓ��D�l�����!��7��ի��X>�ö�w�&9�*��ك�`��t�܈=���{���~y�ƉTX����U���I�1ڋL�֠�<<�s��!u�=?"q�ɬM��n�S�ӣ27%T�WiqV�pZ�}�����x�BSZ��Uӱ��7�_�Sw�tJ���1�ΰɳ�/+,��
+e	g���+����?��t0�/.˂0gdl`�X�Gv��/e�D�W���L�@ )1���[3!��)�@�{P����~���zp?���EQ���U��nh|���'C�ElM��p�-�e�oW�-�l-��Tuo~d�UY���G�+�{�+u1���99�b^�d���� �<C���I��&��<|~�/їM︥��-]�Fo�΀?�u5��T�T4���W�V�v.�Ϛ�{_8ޣf�p�Z���u5y�o��p���ua�k�@�RW9^l�lNI��z_1�U��y�����l���S}�y�����Ǚ"�RV���~^v�N,�ea��J�T�44���q/I�B���YG�����(�L�O��ӿ�����q�H�0X�Ж058i�eY�s{^���z*����*���u�"dRWS�-Wi���l�־�͢�൪��ӵ�RB��9���5jI�)��6]��؉Y��̅�9��J8��-ǲ�bP�Z�S��t��ө�w֥�x�tUsJ��}��g��D!��֛��Φ�g�EU����V�
[�\��5�=@T"����v]B᎖�o��4����y�b,�����̟��e�*N�6��1��=�-�@�(L���o�69�[]-�(w�����N�gզ������6��ҙ��F,7-zWZ�X�7��K4�4]�q?�D�e�[^�F���#�ݖZ5���������x;�o���|�:5/�(������sڈ!׹���y��p���Js���,��Ğ��,�]Qf�.U!��[�=I�-��~ �.'h2GW��4z���������"C����7���	�/	���]q�[hqA�~=�'ft�T�R*�G�G���ϰ�/��nt���V�q��U_eԆ=HH��J(k����6��fO����������kj��0��oSvc7�e�����=������K�<����u]�y��_�lz�\���E���}��]�=�-�����\�d^LL1��LW�Fy�[��6{�:W��b3m��c5�ұ�Ǹ/�l�~�DCgԥ/��u7o��=ڕ����<�U�k����*N�4�斫���,lZҳ.S5P�d�y
����S$�{c���l�9�6���z�K�T^�����[س�-���z��X��+mh<�A��ؽE�X@LvPv�N?��4tEr�{�����M_�����޹�W~�Z��%gN�{��[���R���Ub�bcv7��T�5<� ��v��u7*��!#��LU�Ko;8#�;������}n(�:��
W�-���WY0�߅"�_�՞'�ߏ-+��to����G�}��uN߻ؒ	�{�?�t����Gjo4,X͝�˶RuTK>iJcUUEmD�d8����ت���s�
��Ͷ���.�6c�2���Q�X"�'�hM���Y	��N�@6L��d�����l�p��Jg�LD�����4�g�#���H��p� �x��u����X�x ��i��6��4���:6�+\���	��S��7��E���1��N�fY� �(t;C:�]���%��+7pIftJ/�§S���Zz�"π�es�M?Z��h6��E%�l��ju�����X1�5MJ�7g�}Sި<^W9T����2�%�̖@CD�����\C�k��J܄���#��,�$�L�����չ���ѭT��&��dL}���0ř����;�%�,��C����8ְ�;OS ݛC��U��EaY�8���Neĕ~�E<��1Vn@tʞZ�k��,�	
`��\|� ��R#K7Kfs��(�-xk�]Y17_�>Ӑx�$�M�%ݳ��~�4������Tg��9vP�J��݇q<}
�9 �6)�l�r��,��'V���Jж/�p:�P��g���S�GA���?�Y��Q-g(���t+y��Vq�t#��:ٜ��Б�8}�G��Wڀb@7����� ��t�N�u�����F�_���pIܪ�{M�ci]ױy�2%��g�F�Q���K���W��#���6��ϟ��Q�Cw�V���6l��a�1f``;���߿SN�ܶ�EK����}�D�ĭ��9���h#9�A:=���s)'oM���g;ozy������"茭���M�aMMj�]�&�&�[8��`9�D+�������i�#u�	QҨ������Gج\� #�L$d�`�e�\�Fv �п�����$Hm_��n�+�}V�_9/?�Mǣ�f$�����)�4]�����vJJ�|�
wUVЭ����,Q<�4�*�o�X�IGm����	L�|��M����2�������׆��Ko��cw��u4�-p�����f�����/.YKC�9�6,�5���cL�{�ZE !��ܒ����sˢ��|7�÷��2��w2����ǡ�ԅ�,>�E,�y��,�-=4��VȜ���$6XC��2<��7s�{�Ͻ�ڳ:,�u� ��Y�8����dZz�՗�~u^[}h�FZ��P�YK��@� hz�qOY�i\X���a9E�G�|�WD��%zY�������Y��C����U�`mIضװ]y�`�P_�TI­��ś�Tp��g�ǅ�=��m��5F��z�U���5�v�����7���7��B�v�ˍjRT��^�H��H
������r���*}�l�B 7w�TH��US�Ɂ������O���!�����:M�2,,�l�����sA'�lL�J��K1엠��L�������i��d�)n!8c�U���kC�v��������E>� K�����nb!0 ���%&�#n���\��_��k�z�|��jO=z��B�������hߒ��8~�uc���o�9H)A�[LVƆ�qx����8mO�՜��Ə(f��@�[��Ss��l ٰ���L^�E;����o��AJ�77{9\\1���7��ф(�q��h6�)���G��{��nQ�����jK�e����o�}� �G��x�v��E�|��C�{u�W��F-��N-�}vàM�/ ͷ
��8h]�8�u�,FGOwqyGk�8/�����	Я7A���I��F,����60:i�>��H��&븼��?\����.�(��3�鍬�D�]H�����αSន��ݣ@���������vW=�O΅����|Ƿ�b��bj�Z=�nH���~�;���/�:��:W�u��jm���� ��N��������9�d��u�i$��8�A�Z�YF�{,Sn���\y��CvB��,�j�r�w�Q���r�'U/[��=219����<������e۶�jPa�p��Y� ��Ȓ�J�I�d|��_�h�����s�e��Χz���6c��, 6�ټl=eP?����m�8yK#�h��VnBBK?��&_��R�d��'B�U���eO,��奈 �5c�/N��ϊ�<a���K�q��zD���Y�T��مt�3p�N���0%ھ������KE��[���t50ETYX8�Xk��HxQ�K@��%\�����$���
Z�O*��ZyK?�/��1F�ĩѥQ
�
�mx��4�׾D�ak��voc��3�=���.W]_x񓁍O2������}֙hH��e�`�0ɔ���"藁�h_����m��Z@�K���d&�D�M	
�-�K��gk
M�R+��0��|����*�Ǔ�*��W����V��P�;�2��6��!����t\z2œ8=��# z�~�'~����:�]`������V>+��5�N����0*Q���j
��M�D�q����R�����3\��)0�B�D��R2]�w�Po([7�1O����/O��ʞYY�6�<R�@zK�Z�Q'�u@��^4�%����� �5R
�_���u����銝��	�-��u���~D�tû�$�)^A��;3�����Fâ��G{|;�:��_o��;�p1����X-���C�&&�yq�fT�Q�kT��D���g�:h&u*.���ݕ���b|a��n�a�4�:19\�ul�3FvC�N�c�n�r��;6���mK7��*�� P�݈�g��b�
�p-Z��`/nG��5��`�>��U��y=��c�ܢe��������v1�����8�qD���*���5TMsp��E�#�m�C�-�a5�s�A%M]i&�����J{���S�	+�!��`�	i7���� �'����O7 U��u�7)^����̉3�e
"K���UeA_v��kL�-:l������u��]����K�����+�IH;D�X.�#󠳼M����{�)~��	��ɨ�(1|C�t%1��9��p��E�z�xҠ` �>�5�ض�Ks��t<;%J�����颇e:�/�K��u?<g�+�$�%�Bb|Mz&~���ox��5�����N��>�p��uV�)1ҫHR�'�s�G�7G�%=�\����W�=����à�4�|���ǯ
n�:z�b4�gT~ǃ��C�'xQ��6Ug"T�w��X
����m�=�xٙ\W�~�#]n��aqd@�HpC<Ɍ��w�61\b>��x��
�OwvY'E)���w��G��ߔ���\�v�M?*x���H�q���B��˷�C�qf��+�F ��o���2�l�wO 0A�k��q|�ƹ����yC ��ng_�pc��tk������r�HI�x$kkqo�9<u�8F������}�+�����4T.����"y�O*m��>�`������Yo��}���f��gf��|��c������k��Me�:"?|�U{9�BM��y��x��ǥe[�ڿ=��x�Xn�*�����Ű~��$,��=M�)S�.�=�#�����M��� �)�	�$���3��tnf1�PֺJ
� W���W��>l�d����N�v	�#y��Qf���Ż{�X]��Z������N@PQ%]�(l]tZ�z�7۫�ʪg��f��Xd)�:Q�[��.�"v�cө��($E��rt��MY-�G t��M�|w#B�H�_�aF�;��}����C���K�d ��7 ��E¿�*����M����9�tI~s�7!������4)��������hHc/���x�e��E�%5ز�k{H�ի��o�X������>�r|�
�D�ݽ&QA��rly�B�������9�?�?7�t��+<���^��l	mY��R�W�Q��S��'�_)	P�)f�o���3���ȗ���ʣ��}@,^�"�R��휈�����ZLU�D4�B��9$����lrwD]6�L9��B��V��y<�-6*k]�"v�?��`�t�-�v_{)MD��~��*�{-&��=�u���Ѫ�Mr^�  �ϑ�������N]�9��iY���릨�Lv��M�`��'�K蝾�&��V��]��3�}̗�����٘.(�L���VJ�>+�Y�]��6|�+fx�B_V����X����TO/�S`$�w�=쓜�I�x@pr·�*��E!Q!������Ea1����]��Rs�Lf����g��l�uj��@s�15Z�G��v),9O��Е�v�7FD�Ѻ�9�:rz
�ҵ�����>���;�EM�Ḭ�?<��-�}��ϯ�p��M\�4�y�+�m�S�Oa�v���@�Ĵi��K r�U����9h�xЦ��%�������G������$��~��j��99����L �H����M�#����|Y�w��om��\�]�z�_���WBjbI�Z��6	��lf��Q�s}��k�L�v"Հ�yZZ�M�SUu
���N�Ə��Q�e��yD4���tz\��)\`/�	Ïh(���6Z��җYXX
 �Sݾ;n��e���d�7vc��ꪺ��^�y%����#���j��qtEf���	�QX���&�����A���^gӀ@9��mO���.E�Whhh
����H=R�����S�)����	"#?t�o�a��ǵu��>\�����D[�	���1�u�Je���Ri�e+>��I�[�8W�E6*j�M7�����4T����9K�Q<_N�Wn�������Z�&�2G94���5Qb���Aӷs���ǟ�9����r@`�ѐ.m�B<l �&��<����e�ӕ���C� �ܯ�A_�D	����!*W�!�y�Y��z����ґUc�g�K��o�^�GVE�Qt����� �m�3s��_Y�/�"��#���n�M�~D�{�h�ZQWv<i�V��F	��(aX����XQ;�ω˥��T���zTbrj��K�+�c����9�&/��);񒞡����ah�Ɇ�3����^Jy���Z�5��`1�|& "w�Apk����Ջ�$�x]O�='��ӳ��~�|�C�ϼ�J{����A�����QǙ�ͤ[�(�/%��=i��.$���V���d�e��?"�����6֣2/�S
�@>$����Ӥ��v��릣5�Qz���"�/��`�F�w�g7Ct<�X�o�N^� L��Uj�:�9P:����Y|��Yg���U@�c:[Y�ɼ:%�whؿ�����95<z�f���̣r��מ��_��m�")���b�7R��_w䧜�k��ꆜ�9U�xKz`�gL�����M �w��u�<x��BHG�/��-����"�65o�rm�����GF��"�O���F��"Ve]�5�u�ę%o�c	�C��S�#��T�|�-�ud�4zlW���І�4�)�^X�?C�,ؚd���(F��d)�Er��>�����?��Y'��g����5י�T�+�EI��<���;�P�\G��,y|E��;w�MY�jjU j��eDl �]�="�eU�;�z~�6??���?6�x�d�V���9s��
6��d ��&QQ
��0o�f`��uyy�{a������qa�k�+E>w� �?r� N�t��4��vQ�&;�5oO�#~(Mp2�!hI�ۻ?��$��n��xz�����s�ő
a����,
���B_s�}��:Rc��=�/oT��}&�&8% 4C�s�B���q�����n��Ko9�@	����[ݲ��XUUϱ��.�����-����JC�ӱLA�'��PJ��������h&�Xf�ZP�b���� K�hZ��iF��[3l������#��Eg<г�;]��:�*�Q��a_H�#�C���jgj����I˜̢T�:�O���H��f�zjGg^�����sЮ5�na������.\Α�P� 1'}���=��0�����d��e� �Ι���<x샵�z��⋄'�,7��F[�� P�w��s���y`^A.������\n������gI=Ed�4ح�_���o�P�4��%|�4��Sx��}�vk.:�0:���}�5�u��~ �7I���I���h����`�I��l�S����dK'�.�e�d��-.�fQ�J�;\}d�ж���H6����|����3�9�?66�#��_:��}�prduj�#���h/:��3������pP�^��쒳��-�-o�p���%���؟����h-��ۨ��:��������{'3|�U��������H��3�M"�'�Q���_��Ҭ)������̻{����uu�ҋR8NU�0`�����@"-�I>1:r�2�t��wa��-_v_J�%��_�|\�J�N��y�����a�p��6ٚ�MY���;�����w���ق�����x#�����f�1�ģ�E��^�,��D���9�i��]S�����s�����ի@i�Й��<�2[�ה�s˚i죨xOr|��n �����?/��>v��x�ÇR�c9�����53\�#偹!���W�E���Tjl{��<g8��T��ʾT?~U���(rM�{o��/�e��\�:�ψt��7�&9��o���pŐ��B����2���Ֆ�u�T��w����/1瞞G���e�������M���:(OX�HiS��K����j1�;�����~NT�ո�p�5H��vX%��M�0��8l݃�LѼ"��]rW��oq�#�9%B�蕞]��01A���)���R��j��4D�K��������c�e�}&K����p��{Ç�����dG��V��Tyd0��J���Db�+g�����͠�|\9�I�^���\-Pg8���9<9�0脬d}�1b�o�6֤��4CL��0�����-�!ӥ�l8��M��>�_�>8Y�A+��f+hYSZ��4"�[�>t/�*�d��?B��Օ����?^k�ĚT�y�B9o�������.!�F������<<�=]������{Lc�MC���8SF����������[�^-ܵ��Zd�0�W ��R鿏qoWV��Q�1'e��*��~�o&\�����b�v�!��;�ي���X���θ�2�)V��K��T�>�kg�d�cL�h����,���P2�w4�-YX|z��Ľ��$�F8�mkc7�k�Up\Wj�[�{B�,��������Z-9�qF�T�B�J���ͥM���&&�	��)1۪��j��<2񙀿�>X^j=~ˠ)��b�c �W���a�� b��a��3չ$K����!���' +}�2�fR��Y��d�28�� �bd�X�3L��
��Յn�S���&�Qc��Y�c�Sཙ��i���Z��[�)O<Q�y2�d:�̌�	��-{{�kK�g�����-1s5&<�t���*�҄�����&�xĳ�35�٧x')Y�z|aav�b��(yX�;���`�^�g��v����HI���z��4M����X:�:��M��ϛ����1'�v��ѥ���.eVRO2e���5f�S�vVo��mG=���Gͽ\����3I���n�B�-�8����l�O��dPfه"�m��}ߜ�F�<[�����7"[G�hr��:\��KtePt��YM�����uk�ÿ�Ì�Z����)Ɣ���Mc��r��4��qZ����$`����,?5Mp�Am�m��<7x��.�Cf�9����u��ODIɽ�9ŕl7��1ѡ�;X�s�
���c7�zek�4q|��i���ݘ�?�dq�6ظ0q�L�ah0�����`��/qY@*��m�$W�OY��ԈW+u�s���|<M2H�,_e��ڥ�d��`f�-��O�5N5/��YE�,H� D�&	]�����:�qY蒤���ڈ�ѫ
��|��
�3���(�Ϯ����.8%p1Q/[!Q19��q�Kp�:,)It���MW9p��I���LD��%���"nC��չ�8s|h_3���l��p�ր����_��;��7�t�*9��0hV�i�dO����5�c�3���xޒ��Z\i��&%ӫ��L	k�e�����N	!�ʭ3�:�-y�2�I[���`��fdB��Qv����N�A�sY��u����_��;h��(�R<BIޝ���l�d]i�.�I�e�ʝ�mԷ�oM0��1ŗ�_�fA�"sZ�_�����<����Z���6W���h`��	ɟ�I����j���
����]俶R�4P���$�L�,�UX>y�UὪi��M0%�:+#;�z}���0v@�ʴv��U(�2����H��G_Q�(Dru�%�4�	�@}�����_�kk�=RP]�:�����}UgplU�7Y?T�98`�1� N��+aj��Rii%�(���.��Q�ה#�/j�-��6��((��JN��-��������sqǚ�M���c�N���xnۗ)�(�tO��nI'�8`k�g��r�.."N�@���� ���_JJ����~\�z`�L�&x�CM��s���{�9b�������U��U�s%ܳ����a����IU='�:�:��l�`�<�� Vz��?1S�Ygc;���0v�˓�?MJW�_�>�V!)Y �X-�'���C�_�l	�I���ܿY��z�N�,c���.?��6�4G��Yc���K7�=��D6K��)r��"�OJHGP�=��K�� ���y��QѹZ�q�Z���515��+*�#���[b��Y�e$�����3�j:�8�-�n��)Dꜘ�6��:�����==`O�~mFP<uAƷ��(��j����0U�W�����'����\��]��+s�{�3q��d9�(F���z���P`?�y�Q.w��##�VyU����rCWL_�;\ ;���@v�P��L�,��vR(-�N���A�Y���I�ڦ�(1Ô�xPP����h>���d�e�H-a�օ�����FLB9������q��H�|�����W9%z�?@�*����QOV@ൔ��`K�K����f4L��� 3h�NM��'qɛ��QC�n�������+O;/জ�eS�y���m�<A�;�%�ǋmCq`Dy��7z+�/#��w��Რp�/����q�c����$[
�u��Ϙp��<^C[A�@M��U�4r&Yq.�x��7V9Ƌ�is�ma�;�� ��2)�^�����4$��<3��`��;}�DZm)^��|�Ti��YqY���j�!�*���2j����ԏi߯���<�c�v:�s��3S��>�Q9�_Cx�V�����
H�z�-PD����K{�ӝlZ\ARF@�*��](�'K�q��'w!��g�����~�u4A�{�ܚԂ
"�I]��8	LR�����k�P�s�u�|JK��n�;�1�)'EF`�|��K�.q.��H�_O�p����C�ꍗ�-�/��~���
wNw�� Τe$���a�A��<�IJ���[aw
��S5U�4U}�M�����v���_Exw K�b�l<v�0�fI���͇�aT՟�2KW��S�j��c;�dK�#�Ӄ+u-&k٠4SS�F))��wl�SG�8��Ő�}Ͽ-\��tB�)4����n�����'	\��65�ůM���מ�y�(��y�Q�(�۝(YY+oц'S�f�����G��;A�'��g��Hq#8w��Ȓ%+��4%!A��2s�m�o�Hi�I���8z�18`f�d=A�P?�-s�A�ϸ���t���;�Zf��D?bx��0�;���JbRxP?�Zh�_����K[.��&�mp�~��(����C7$�W����D���8�}>�hn�R���k��Tf�M�^S���D�+&'�L�x�%�|{����n��ʴ|fE�"��II�����������e��cC�kn4	��G��g��%�>��N �~^���kd�x�Z�d��"���^Q)���@����s������� v��/��h�m[8O�@4(��u�HME���"܄E*�;�e4z��=B�[��w2��	�N��D�C�Qk��_�@�����y�::�R�ܖ�:6�4��r�K؄K��WB��J�8|��n����Y7�����a��mB
m�{#;�#_X�s\o�����nt��x��׏����{�C�O����T��m��e�/�Zk	�5�[�|z�Fq!\�<��y�}~g��9�GB������N��0��ޡ+�&p�D*��-��n���E(X�lۛ�>�.ґ�X>࿑rk��������/����HI��d�u�Խ��� QcI�Rg0��Q!�Wsq{�O�4�vԕ�Wc@A�κ91j�^jj���חB��D��E!���?��x�K��	�N���k��
?�c~�=���D���U��!�Ң�^R�6m {j�W��5	�er����a�mu�z�b�lS9���ǎK�<�@C=�4��в4�����ԏ�T�N 1+#7�6R՗Y4��؆=^�"�*HW�>�<�{;Z��lbRҿ���k'�#cs�rm�y�܆�l�A�Y�b*��y5�q'��C�2gc���ѻ��lE�r	G����~ycҧ�51�@�Z��6��.jL�nԜ:��_�-�u�Y��z�?>�V�B4�U��||Z��~�����{PV49 �9�z3�c�j�Ƌ�R����̈́�d{$О��C��b��%���[��I�}UC}3�Z��j}��di���	TX�ʉ�%�5��T*(�Q,<1�H�{��vyw�^���&y���"V�#�?P��r�/D"!2?ޣ�W���ƾD^8�Ys��?b���C�3���+��h1)��c��n�A!���W�(=XU�8�w�.��du�!@/
���;y��W|�GYؕ���i �>7>��pj���������-u���g'�x�!<�x��x���,+��50?M��'S�t����]��>��� �
ԈГGhȨ���D[�I���B5&�N����E����	@��@EG �����l�k�������D3B��W�׹�&�p�d5X�S�.#�ƍ#�5+���x�L��<K<܇�F%�P*΍S���1��0���VGk(��Ӱ~v�Һ:5��u�r�ܬ�I@��O����R�n%����~�Ɉ��d�M���I��v.|�W���'�UN�.�=uk���x(>,c�g�H�Cw��D3i��q �3}�J�8�>x�=@��w����4�Tb�v/�*�X��x��K�����5��I�����8��n?�k��'����u#-� )��%9Q�6k�&��41���[��d��<,�\�����i}�Zcȉ��#jur���_�(��^�t���o�g������_¼S��
�<..6q�-�j"JI}F�������{ao�|ﳃ4�n���ԣ���v����T�^�9�o���^�tI�p��:?���H7v..��\���$'�.w0��?f*J�qv�!��%W�l��cue~�U �u�N�n+��8�(Ek$ob�OF���P]�����;�]3"�o���*+����c��5�������\U9Vި\�NA%#;.,�3��ਏHo�;=Rt�H�/q���<i��K��:~!��":J���j��/��=���}T/���{ϥל��2 �p�r�|K��UP�#��Z���ZWzSn�Nm�`��+���}��=�N�s��3�҂��#�����$�������5�Nb8�TVE)�=�Q����-����U��4I���ſY�0ƊW0��>�O~��&l�W�äg�/q�S1#���=Y?<|��,����'z}T�G��X0���8q`*-����_�5Y��v�x���>�&z�G�u;��37�2&1l�P���䈌�,�|�0t{H�P�� �6ش\��{G�i�a����a��j�2��8N\ ��y�\�ȎF�&�'~��E��e
���q\��K �U=�t����Ĥ��&�"L�1>��s�%Y���z!,9�k������w�v������4��;�˻|"Bv�v�� �j����$�y?�'N�j;EN�0cb�_�0����J���C�2�����̹���w��� 7	�π�w���D�M�r{�{{�e��eK�2�>��v7��G"@�����=i�������¡/`�.��rl!N��j��XB��K�G궪Aed��Aa%�����9t��Vb��d�̠z�P���PO���P���'� �RyX�dō�E�?P����o��O`U? w��aU���y�M�њѹ��m�b����q�3H�)��7����Y%��.ƿD�_"ɗ��/���J>с���D�i0���vť�W�J�|��y3p�`�K�#y9#ԯ�D���(�l�y�Q�[�L��Y���{`z���ԗ9\i���Iw����#0�-�iq�2=���B�8��l*�l�9�[ �(��ϔ��ՎK���x\��Wu� �_M=+p��8����У�ɥN��k�I��P���Pk��G�&�W�����b�%��>�G���s������*J�)�=	'�"���^Y1䯌��P���IĈR���-A�d�:��Z_?P*���}1h!'����9�f~c��>]���"�S#Q��f!��2+7�
'�nX��	�l�5���As��|�qj~�LDt(�����U��K���b?��S�4��Y���e�P��n���AP��d-��Ey`�*�7Ӫ�j�Ƃʳ�����+��SV��B�
�@!�.q^�9=F�ݛF~prZ�癊RQ��R���77���h�W
U5搿���Aӊ��:��<Пj��L�s���I�l8���J;���#և�J-�Ӟ��
W�0T�q&��}�� �������Xw1��9U[ӕ{��\�tt�p?;�����0���T����+�-��Ǐ@Ux#/O�Kf�5�����w^p�e��7��m��.�}�&�߭r,��1z(���F�-��r(P�|�U�q�y�;2�=�N�����}݇�ؙQ^�ݵ�f�L�'��w�kۑ�**o�����e����1�{i�d��􅖲�#�l?�^�� ��6�+�ti������A�c_ϑS͛�7��rtk�#Y���\����p��t���H�
�h��KHH�����ㅌw'[���Ό�q_z����.�B^�ex��h����u�	�f�����G�����T-���Y�X�\��#(�1�jh��������5���yjC�
=f�s|5�%B*��νei��G��{���ݕ��W2��Ծ��㎿0��l�ڷ�p��������\���<�Wa�P�Ym����LrKl��x��P���ˣ�<���dmC�v�9&���uиՆ���L�5���ܿ�e�F�����+���������ir��s�3����
+?J�^������3��2�(� 4�r��'��J��o�uj�	K���w�4j�XD?�ዂ܌p}b�堅��W��
b�5ߋ�u��W�֭�g�&³�.�v�����m����������8�R�.w��X����t�Z(\�/�NL\�Gy��w��C.�B��;�`T".e�\�\�+��sK�'�I�T��<�k�:��� S�����&�%���-�)|B�,C��z�!��2agU^�����&/���~�.\|V;��Z���4���lY��qJ����J��Go�m�'��WD�.�&���1~,1R�u ��h�*����sGjz�R�b�s]Ӹ��.�	U�V��T����ϯ�6�_�PV�팶>���C�ۼ�'K۠�;uyo��OX�'[�e�48�Ų�BMRM��k||������o���y\�{���W������<�<>U�����f�1��N]�b.���3*ܭ�x���$��nP��Xޘ��]�ٶ��sGEF�׎���J�&Ql�C)ܧJU�9�[>����-J�%-k���y�0jbb�[����ձ�Unڨ~�㓡��S��d!��We.���N�T�PȮ;���y�L��׎����-�p��B��`�{~x~b �ƅ��R�s�M��	�G����֞�����
���a�"�}Ibk��n�f�����3_�J��r>{��V��l��*�8�aI�t�(��ym�u{J������$�trE<l��٤"�:^�닕�/�),��WL�8���LQ��
��]n��:!��z�M~o����K�����-o�\Y���{vJ�>���}In����p�x|��o��[͟N��[��{�89��f<��̓���e���
 ��G��7����4�F�W���\��琁|�F�6<6�H��Ր�U5�v�+�}���޻�
n(�\��[䢅铨���Iz���.���sYy k�Q�ܓ��ʕ���1Ub��po��o���}�X�k�E-/vv-���n����͸�eKD��r9֚��|0}��k>����آ��� �X��Zӹk��K�`0�c�V�-%6̎ƒFjK&Z/�аH+Iic�ߋ�N����[/���^e������&�2��Rծ�5�Čq�}�ƨ�5yGv'�8V��d�8�������!=��"6� H���o��jg�U��t��ז7;B)��(�Z��l��cO��ʋ=�	���fR%XB3����E��t�Ƀk	=}��a�-�+�>�7���JJ�P\_�ӵ[I���idpn9���n���#�a+��;+�������×0A�I�U&Jؽ��٢�o�q�����}���&�S5��v�Z̵�[b>�zn���o�p$�
ﷆ�>XӚp�{G;o�-ﲙ���@g�fF�`3��Ux��CO�W���p�Λ��D��p�?/1�nSO����;�`��w�߾�8,*&�l/�.���=���߹!]CKA��;ò�pS�K
�pkKN���3�����/|�[[��&�/��j�xc�3������OL�Ց�L�O���0��{bl��U��Z����X��P�Жr1�Ǥ9HްǸ��t��6��j>�^�_���LL<~��3�	R�h���.U~�K�=��l-����A�ՠ�?�׿uͼ��[M��ߓ�^nm'>Za��~U]��=<�PhX�i^� �%C+�>�n��6E$O�vfd\�L�	ˮO'.*�ºDdPۇ�.[��쯿�̿�x�e���gN -����kM�{��~zXޥ,Yc%��if䉡��]F�
V�(
�!^ǾP�rr��[�_ V���G�vv���ݗ�!j*zV�9�UL.m�OV��)��*p����fw�Vy²L�k�9a铠Nx�Ldurjx����y>Vh&�B�CO���L�g��s����kW���&l�Ѽ[��j�03�4��%5siΟu�<�b��X���F�����t�wN]�	9�{���&�!���t�
T��C�C�[��W��_^���<|a����7��7��O�Rz{~�$���Zx���ʙ*;ȩF'��h��6�R+��>;5q�ݻ<W�Xc����o�?҆��)�C�Q�ys���J����m�m�E��]��������7��Q�b.B���mHMH��8���b�@�����?i�O�FB������o��[��r�4?ㅴW�����9G�93���\���*TT�Q��</$(��x�-3^��"�G?�G$�}���˖%��n�$[^P������o)*�o�Y�j�p�6�:��*>n���_���F�o4!�)L�D|���
f�0�J�>.����fO�F�$�Fs��䆆w|����׷���7�0��K�P_�&�Y�F�-n����S��+t�%��>I+N�s�iN�������Rn��#��0.}�l1����ci�ͣYv�����H���.f,�)ĦDP�>�N�X��_'���X�bF��}��>n���^��ouz�/���U����ƽH��Q�G�X�M��-j��� "���k�I߃�Ȯ�x���:Z��ճ�xq��[���q����{/� ��5J�����R0�<H�2�Tk8�͉��?mTЮ��:�l~����N6�ds�-�ƭ	�3%ne���;Kϸ��/��,���
,I_�Y�e�؞��ga�!��� �����(}b3q���� ��(���|��W�$�o��=GR�,����3gߓ���?6�s�S;9�3Y�����{?2
AԠ����7��9R^��/���U+tv�.�AAȸ���L�ٯ�)�I��i��M]E��U)o[ m�9>>D 5���N�2�	�'?�	fE����;�C|P�I~[s���@���Gp�NB��qm�m��T3��D��B�}��\j2L�b��e~�#�̕t�+�z��6;�M�~�Ǜ�~��\�?���D����@����?$30�?\�uTT��>NJ	8�J�Т�t(! �  ��C���(]�tw�H��0�4C7�;�z���}�õ.��s�����~��3(�Y_o�=�{�p;�U1���Ю��������_������Ɇ_q�װ��y�2�`����{���w=|�S~� �UxoOa�9�8?
�E���5���3�cUq\���Xf���`D���~��������#�k'���[�'�Mg���R�I7�`�7g���N�5<�v��*��I��&�G�h=e�<��}�=���fo�m�Ԣ��2\��y¾�A�}c䪭 9�x�"uR��)a;dnj�d1ht�񾙖�.U���{�OOOb������>�Z@�;�w��bá6�{6�r�w�kng��a4�G���O��z^ 9��k0��t@W���H}����\� PXmjMC}�x1�E)z8��C�����}A�������6@^FK���n 0Խ�v���ȹ,���muP{��e�w��zt����F�����-��iap�8�>*B埒H�_z�k�.���*PXc�ߗ�YQ�8�������#�a���`��Y�x��2��mx/������p�}�gD�+�L'�[�&��#�^��R�ԸU��6�H�婷rmE���Q=�=�)�ɑ/��k6-%݋n_֭$N��� ��%yc���U��p�n�A������s��v�Sm��_aa�7�O�`�Hl݀t.�e)���y���+޲_�m�z�p������2�����j5;q�|��`�7cG��^�����r笙�n�b�[��>�V���ɻ�%�ˬW��.K!e�sN����O\Ra��Ig��lg�u[6�,i$P�O$!%�q|��K�4ھ>�o'r�s�)�����U�NЄL"--Y��@������E�4�&��YX{�w����.]�Pۥ�F eM*��;�ifR���Q�;��<�?���X���@�s=ʂI�`���� u�ےp�_h,/�R��c���I�/�R ة�~���а/Uw6��"����=�0�Y��rm�w���:��_R�CL��!�@[���k$�:��������I�4Zw��.�Q|c5$:\�%�W�@������C�%N;��B>�%�&J��8Uw���yقrM^c0%��#�������M�����Ҽ 9��t��/bD��\��"���0��o9�EP�w����dθ��!��J�旉�]����LQ�.��m�@]9s��y~��j��
6x���>P
6I`�Y�}��U�)�;r�r�1Z�VdոB���xL0�@�اa�������Q�q'� ����|>пj�VYʡ.3ˉ%Z��W�&�츰X��ju�٭j>o��d���N��p�fzlUw��j�u�s�����Y_�����sy�:���g��܃�|c���H}�c�E]��<7 3��FY!D���RZ!�`��g�<��F0%7	�p;��|~���.i�K4��~I0�h���z�>P��)�3�,��	%�j�^�k�>�ţ���TV��������"��,�����5�S��8���Kgu\0���
:��0��kQ%�� �=�2p���O�����M�F����؞Z"?���Nr:���!�j�_@@��uo�t�痪���x�%����.	�p���3ϲo����Wfñ̰G���;��lN^��!�a������k�~�)��3;2�4XZpN)������~��ǧ�N����B�����o�k�<{^X�(���(X�@�bu�{B�}����/�,�)EUFMU9��Y�u�@ܻ���<��%��O%�<�5%�"v>G%��XWLEu&y�V��ܗ����{U�T�ZGX5|���4��f'��q�	�!a�$bb�P�r4�
y���G�����FQ�����IzÜ�o�!GB]l���8�_����H��2L'O�����q�D����xg������\��tԯ�C�X,9{�U���}����d#V����ۀ
�V9��\�s���)S�?<,��yQ.�A�!	xq�6d*�*1����	��ad���>�Bl��y����?��:�&�#7�1�[��u�:EMUU=��b��n�
�W���v;�(�����\}_��b� ��w���u�������т�3x�K��z��=�g�翿�D��V����E	(�ߴ��Xq�e���1Yc�F����Ņ�v�:^"�ܱ���H�Ro��=<�����S���������YނF��t�A%Q�LS)|TޓL���t2�4��쎢}p��DA5;{��0+�h=-Nb�>��o���-U"噡�}3��0�ER%E���s���񣬇~�g�3�����G�yv��j�����ai'��]�@�kQ_\Lǩ�FK��?���؃�xV3I'p.e�p�\߳g���q��ȸc12��-�`?�?ɸ���b�°��{�\*��3�5�f{�A�O���mAߢ�y�v*���|�.�rr�\|�s�.P��[L�T�S(H����BGSFmX�5�YC�����·a~ ��gj��LU����*�]1]j_��y
��pݱB�I�S�קJ��[��d��X��|�s�0��W�!,n.��Ma�Iglɉ27����~l�f���Ų�$�k^���?.C�����L�l�p6���L���6S=�D�Q��[��oY��߿�8hZ���1J'yإ���Y^y���	;��f;f�Y���3m�-�t�D@,���m��%KԮ�wv6 $��u�'�U�3>���,�ߵ>�7kp�q�Z:����s��2$���i�:����&����b���
^��hg$4>��p�1�c5E��n�0�c
tI5
ʅZҷ(n˨��L!b�t���fe�3�p������@
J�,��;
�@����y�#��ޡ����ŋXd�=��Mv�e�����6<Tā9�4AVo�Ȝ;����ܻ���pf�b�P�;{-��؉J���B`���`�.��T�{�+t>��%������	��/�m>�#�f�HɨM��8uQ"{�`�2 �&�@�.xm<.~�`��Γ��|��Z�'�0y���
V"#36G�h�|��ފ��o0$F��_��HX�۷�A�M�E2�|&�:	��A]-Q&�jTV�-����8Ն��[�H^EZ(���$J�f���dK;����I�4�G�L�(�}�h��7 d�
K��Ų�L̩]Ϲ���	������k��6ŧ��0=Os!)��t���_
N�3m?�*ΊF4���d+�1'��G6ë��6Y�8����'��v�����s�݁n��"f2^���w��etl��][kg�M�>¡�?��ã�Ru2>��nN �)2`�Z�O����4�;d<�`Zׯ�r�+��}i�#��e�M���;s�%�Net�s��g>K�Su&c���jz��<�N�,	�S��W�s��v����E�>��+g��#���>?�U	W=C�G��л�����R>ű]R� iN�M���Cg�I��c�sLe�W83�}`2[Rܿ��[��6��KD=[�JfL���m�e������]p��J/��-f��ws��to�垂��Ò�/Q;3�}��.��ƫ�l�p�/6�E.��_��uʟ��9Lf���郝�\���ݾ��vrh� ��.N��	)�k.���Z��KX7��!]�o����5����K�;�3������E�tJ�a�7�����[�W)�LƶD+�k�M�\'�*�����0�ܜPNp{$7x<3p3��?��Rв�"��V���î��ִn�H�es�T������K�9-���co�zk�sgRa̇jk��)�<�jo���Qǘ�ᖔ�)��T�-6�
i����+���V���J��=<��7��L��ć�,)�������~��m���(�Ǒ��fHJG�P矛�w���; ��ҝ��.!?�U�7s�z������e��J U1?�s�� +Υ�Qd��u|ӼN�)���FRI;M-�����yᕻ�뒌����y����?L���scdţ�h��ki����_�����װ&vÿ���L'��G��}ٛ"fQ=-���媲.��&3�HE�zZ�;,�%��hN���r�1;�S�Յ�ļ��Lg��,]�-K���;�����Z�������0y1��.�c��-�iC�E�2�^]�g�ѐ�`�<x�xS՟�:�b苽��G�;|�pv!���Md1|C���*����� ���9��mq�u訆�-�*���J/fE/���P �_���i#WM�� Yܩ\����tkn��� b���g邎f���R��{ِz��:����+�B��7&��(n7�!Z��f�N60��%h&&`%�exǣ[�ф"JÚ����cA@\�4�4��?�H�`�<��`��h۞sYJq4�E4�;4�)y�=ox��j���Z�i1���w��7�ng��3>���~uP�/��.�ݚYa	�%�]��O���nO�-��R��oy��E )����, �9�a�5v&K����wj�����&���\��M֍o*3�<A���������̸�ԕֵ�EL}6H�hB�ʘL���tn�Gv/8a�)
�!����q�tԬ�z�5܂��m�S�t�+/�V�Z�e̂8B��.W�Pֺ_Ж
�]�����o,���/D]��|��.�Ł�<��s�P������s�<����¢�9Bq�t�	3�*�p���q���}��s�i}��'�m�ߵ轷:�ۀ^����40�����\�rH��A�lzq��������LY"���B�5�߿ٓ�
u��p�z�|U¨2�>�����<�J{���Ӑ�)C�+X�l#��5���YQ���__�$�%�7�S.��~������Ku~u\nړ�;/+s��4���J'�E�Z��ͳ��,ULN�[�cK.�h��
'Xo�Q~�iA��|�1�`O���!9|V��O��YO��I�&+��:�)� |��|��-�{{jLq�䣼���chS�J����Dݕ��A��^S�$P{���w��;�A`2ږ��T�I�g�B��OȘ��QX
���%@�B�6�h�C����|�C���Pܮ��S���GNض�T�U=ph?�6bW'+T����ݤY$2W��"�c�f��#�0+���-,vg{Mi�]��U�_���X�ϤA��J�(���WT��O��x�����"-6Մ�����`p�K�����U��}�z�aH���)]��Ƴ����V�nI��KP�q�����\�fQ �H�X���ީy��FÛ]��,@��S~�h*TlO��#$��Z*�u�]����m�F+�v��Hsț���x��/hH�}���dSw}�̚�C����͙�N��F^X�r��g��ۧ�A�J�������C����q�>D{*SK��R?�S5�;5[E����j�[Lĕ��D�ȴ���(�E�tD�8��N�W_:ϊ���dbc?hz
��{�d�j|1�k��W�Ǎ[�6��(�W���M����Vr��b�\��xzEO��k]E5�[�W�e�H�m��ڊ8���Մ��V�ܢi���ˇ�L�X�4�[��6_Ua������?�)�����b&�OM4���u����>�N��lg��?\m��Ohԩ9=�Ɉ�2�1�ޘ!�%�l�`Q�`%=�i�����8���C��=�+�0�l� J�����Mֳ[�[w��얈�,��O�V"��K��FP�a��	�]�}���ݚ��0��@?���=k덁��6z�OL�R8_��;��*�W�NSIG|<R���T}�ԟ�^�f��x|���%�x�m�hH�X�� ;������b�#���hQNa7;E��2��:������FQ�:����~��}%�S+cogZߪvw`$be�K£��!#�T6q��R�~@�/*�y��j��N94.$n�?����dF�j���,�\��W۩`����aY�2D�p�\��dAg�B=_�I�̈@�l�b+�27�읧����H��Oi˭��� �����/]�Fk �

gp��Y��f�4�� N��~�~|����~����R��ܼ����ޫ�G�yl(�Z\>��S���%	��@í��N��e��-�
�[�.g�aaa83�Q�K�`�B� �BV漉}3�t��xm(���ژL�s�D���ghI�FP��� X?��n�8X���ڧg�/�ڐ?���������14Uxp���,�l��4QuG*^�'�N��[�x&�`�=��b:���L�ߖ�~yŇΉ��֜�3b'��jy;����Sm&`�A�7�y\�W&7T�?O��i�>_7�&~��!i����9��5��z��o�|z�v�V����������ӂb2��k�m���Y��^j��pֹ���ɵ�ÇPS �a8�f
�:�؜T�1
MF4���cz���?Λ�,������D^�T�z��`6��sz�y��%"n���,a�A�F�/ eL�CL�ܼ;�,ˠ��������5�SV*[��Z���.�	��V~��4�5H�~y��c�c�q��(Tc�џ�M����W.��_�;m�@M:���_�}5���G��S{g&@Al�໴�Rx�vll�r��Ly�W���$>Cr�Ȯ4/l(%�:P~P&>�^��=$������RpZKB��&�,�Ŭ��T 5� �M�&�A���r����tc�}4���~��\��(��D��~���+m$���B�A�56h=����{�@��f�֘�^�!�YV�N)TY�
�L���Y?[��w��/��,�Jˎ�Q�$#������LU&�\���th��K^
��p��Z��Ժ�n��+�:X�3+.f��]������#�3��#J�|��	F��C m�e�ܞ�������������'�+X�D:Wef���z�-;p{�S��l��bc^��!s5�wQ=���Xv���[���p�ڥW�I�gm�Dz����,�W���Ze��&�q��}��F�̧z���k�,_g�D܃9��$og�?A��{F�7�ۆ���՘ў�#��]��I��r�B���%抐��_`^�Xs��������6�����Ǚ���q_���6J���L7<H��Q��2��^;�{?�1�ᙁt���M�^�A��_?���r?�M����R�B���.�_�2�������m'��vӏ� (���!�Ž�Tbw�3��;��a��ڙV�y���`	�E�#�%P���9�rZ�eLܮvsNBiH%ﮧ_�,H�ä6tmK�%%4	�v�'_߅�Q�(x%��V��d�}/����0p�׆�
;�_t1�1��(`ڰ3.�2��M���
Jfچ���=@��J,JЧ҅��	\<���r�V����G���%�&�-���vG=�ddj���j��p�.����tFi�S?[[��1��;�!LW����v��Im�zz��)��������?!���� ���M'K3Ϊ�t{���G^�LO&	�*��e��pVY9�� ��P��l�a��:ű}R�J+:,,X��z]�h��>�����ɚ�ռ����50'ׁ��!Iǧ���[N����R�
f:�m�?�pˆk��nç�^�:|�AD�?wl1m^8�_��%w�.B��.��{�"�4�0�"�Rۥ*l��X���	���MS���J��c�9̔Th�n���B�fI0Gi�b}2�A�8Փ%�W��po�������ʴq��S^I��N�R7�a�C�Ĝg��Lc����"���V�yoO�R�A1�i_�����킙D�K���y�}2hZ�IQ�?NN�nrβ��uz䊼K�zY�Qem�;XQ�c(l���gMn��"�u0r(��e�П	�}����[H�oٜ���=tq/�3N G������#lq�H���.? E��>��Dv� ����0��������q��U 7���5
�3����;��z�5���2����]���Hzrx��(���qy;��)�XM��hv�"��`=��')m!)�bm��dZé�QE\��6ތۊk6y%e�G>����ZSS����f�?�h=@��ʚ��a�oޝַ���_D{��V���B��6����.���)#�J]�B�k��
��Y��E�{ �YE�қ;d�yП���D̓K���������M���~�gZ �uF���|����$R��,�����ַr�4W������X;�<@����9u����ȷY�%�1:BS�y�`�8��?�G�>��ʛ�;�B6Z�u�잚H$�UT$O�l֪�� �f�#���[�򋊺㠇�(����9O;�P��KHӰ0�FBB%�D����� U��s���#D��ߗ��w1�;����
��W�.4�7�K�(f8�H�ܿg��裰�s^�!���1�R7�K��s���k+A��k��(:���Dn���9��" \���������/��؈HDY[Ul~�Is�"WH����^���~3���7��]U���@)��BT�*.{�@���蟏5#��1�O6��~׽1e����v�ws��LN"���;�U_�AM0�G��M h��ȴ��],&�뱞E����?_����U�@J��-b�?�T5�����7-����͡g�,\
&�l�C�q&M�wkS�Ø좀���]�RE(�g�0��~Σ�t/AN����ş���yW�������ƴ�*jv�B��۵Y���-OuQw��Bit��u��l�? ��F�-��fOh��q�$�ŭ���RaK�����4���ԉ��*;?�)��y��[;Ñ=���>7��'v��]����A��J�}� �x����X��=t�����nQ�~�]�?7[%����<� �7�����ߖp}TN9ڳ6J|�n��|q���R7�k ְ�������M�:႙SCL������v}�d�k�F�,8��4C�OzKMLn�j��y�����5�v��j��wNL��ީ�����	N��G��o�ZˌsJ�4@�q<��u�
$��VC�	�2 �7��3g����q��Q�C!(�!�fUt/P5-^&<��v�{54s"�O�<į��om�@�v���t]+(���-ۿx����	䏎��HѺ�����''�:�$m(��_4Oz:���%N���K��2�TM�8��9ƾ~�~c�;�p_V�A����.?����(G�S��)��� g�wl��L��������J��[#`�>�pu����T�\K�|K_������x���Yq(I�f��9.�@Wʬzg .v'jm�_�~�u�?��f)�}Fn��oi �h�j���H\���i���R�	�A9e�W�@N-�db쥌ݘ��| P�tُM�|Q�@V�i�5��׮��"�jZ)�{g�Py�p��m���Q-'� �>9Y`+��o�s�vXl�p�O�h�3��E��څ����J�d�Cɍyč�\�@�d��<L@�N�����I�����ݬj����Ӂj�3�G�Z>��˥G�ѻC�o�8�҃@�:����D��@���A�QW=5
[����K9�_��~=����p^�~��*��U����u�]�zw����YfH�f߰O�⿳�d�D���[��xD����DՏLE�����_�{/�дL�B|����3�f���?��d lK\0����B��afx��n�{�=vVP�Y2�a��k�^
1�f������)��=����A�
�N�o�Og)�|�@8�JR~�o��3��z��U��{q��<Y�����')�4���2^�U��G�mp�����"�y���a�;{��	��m�=n}ѻ�P|����l�������ї�?����S��b5�j{PR ��J�&����?c~�E&�+�t�D�-#��nQ�����c��]�р�*@aO��/L�Z��ʒ�oz��J�����( -v�n����̌����E&ZjX�����t볶�kJ�6���&�e�E��x+�~'Ä_h�\���e�,�2�}�~\w�������40.�>����62����˲�����)�Gh�;Qhta��@O-⎪��M8�Q5�;�O:�>���/��1YL>�0�`ԕq�gɨ���t*��J�a����  S҄Ǐk�A��	�ӫ�ōR����=�;��ݚ�;X����*e���R?��>C��D�w<#�R��mȋ残�{x�蔫��Wh�����/f��R�
>��ㇿ�{$�r���[uB�z�f����+��5_1�R7.,o���׸� o����d�cW�П��?�Aշ<��}�:]5֎>3R_���"K���~8ln�l��H��Twc��%�ZM�p{
��(�������^�-�� @\9��_~0�%��|F��q�w�S���E�hհ���M°�~�w�o����(�|��	*W�Fa���x4�
H���_����9Mj�M�%] Z��#��&3����L���H3��������Dq@����i�����}�'n�z�r��9�ݬY������t��t*m^ɧ�B �uKw�8k��|��vF��,*�LXɳ��v��c������^���lO>j�%�{��
ɗ����J��z�v�(r1���lYh�*����w��[���]�3���=՗	a��Yw�C9yjظ�����Nc���N����Z���ט4?�,-]�����3��Z��5�qÿ�N�!�� `�+7�a����ۖ�����V�F��a? �L�V�j���_��X�%L�X����&�����󪱷�/U��q��:�����n.��-]�Q���fE��ȔƃO�7��Z�9~-zz_d���V?rz��R�h�����QP�̻AvhN�X��T!��߯�_����Y�0M��|��3U�}M���)��?[�a���l�:�ux�T�A��%��w�8q,ID��^g��|/nQ5�_�
�3�t�\���9Imp����=2��X9+Ú����w~i󅰱��+[���O��r�4���>V�V̜�*��ޘ��!f�M���*Bm�<�#�>)�L49��8�{�;|Г2�L0���~�I/���M��|l�UU��^u��n:`���_d�z��nws��2��>�����f��x�'�P�qWK���!QՔ��pb�V����h$��ם���N���uF��z��V�S0U���QԮ�jt�S�$�cs~���t��-�3X	��񶥦����R��K���['����3���,!�j�����D}�Ýl1��ڒ-?O��L?G6C��-a7�_	\v`���j}rB����>�,���+Ϊ����~%�k+ ��dH��^������D߹;2�iAE|���۲'�4<X�^�4~(���
{BĊ	4�	:҃�b���Π��%K�/��Ǖ=�ˆ�d����,m��[Z5�6fP2�Ө�א��$��3351�"WvŮg��;%Q�PB�$����I���[�YĤ���.��w^�Ҫ:�<����M�x�jN���^>����̏�0&��@d��W��
O��8��6�iYњ���#� {lv	��]Ϣ��ÿKA��t�8�}5ԙ�د-_��/w&�3"�����.�!P���`)Y�_��1����7�H�l��EԵ=�GY�hRcs]�����ڣ�D�������E-�U��P���J�gױ)���{Ͼ9�����ࣚ�7dl"ɲ}"��5��eF��a)�Z�i����YQ�"F ����{hd���7V����l��Y[9b��S^��%�M�����v��YX�����D���>洢���z
�ad�{띴����)�(��s�]��0N������Ќ���Q�;�,}H죌�Y�#0e�lo����4_����Yc��9��},��/��s=��R����n����-�L���8�s�{�.��1rR��-G�>��nO�����-\	�2u;+=rB֣��l�/t���!��b��������,9v$QPr(��0n��_O ��ںNc� ֺ�v�Ϗ���u��rB�8�����a���A��u�U�T���Ei�7/�6�V?�o(��^�~B
y��߮���� �v�GK��̴�nɵ�.\
�zt8��,����ED�j�v�5�x�w����p�K�h)������QF1���ݷ@�^�h�>�>�#�.qYdA�ry������AʏвM�7^!n�3�u���9EM?C��S��^j(������FGMK��Cj�I+�5�{��v�4�����@0_p̏�Ί�ak�5�Oz���<EÕ�148k�`�6�h�;�B����F=ѣ/sힷ���pW�?dw���l�3�� �%�����-g�v޿��I����p��є]�?$�80:�Nv;�Z��&�L�1��L�V����%#A�˿�5[D����A��h�d��h04���"�����Y�-s��q�3�_��Q�n,~2`���t!`>.�@��l�;w�l ��&�T�}pjl� H��~8��&�����5��
�p!
���~P!�d �0�p0��	_b:�� +�d�s�bA�+�ݠ.)�K����d���_��|��J�LZ�A"��K�]!��P�PoBx�-!B֤Z�}���~��cv�,�����2��#�"���ˑ�� �ߥ!�%u�Z����j�~I����';w����I!�h�> ��}t���� �s���6�:�L�S�@ ����c�F�1��M"A�$�.TC�-@$ce\1��%���@�w��P�M��4�Ŋ��]8�������.`44�#3����L)Rg���� xA
��"ؾ��)'�O�&T�q
�{m ,f����ۍ�Ʋ�)����+��Vѧ`�f7�Z��/�>��|T"FP�D�'�6p�Q�y�]U-`:[{b���L����2��cW�����H����)�
���ۉv
�,�'$`, ����J�ۂ|v,w@HtrbX�� Ͻ�	F?g����|$
`:bR)>F�[�o�1@�HΑ�(����ٻ�{���w9�0�8}pAەόS�`�s�ǈQ����\E}}�՗nn,��Q�4�d�H��g&�-�&|7���y�������e.g0��������m�v����X}� ��@C$ܑT�A�n��C�X����e �H�����IB�~�Һf�n;��"^9�w8��2r��mF{����B����Wݷ�����z�~�w*�'���8�s��3z�{�����ɸ@�CI�R��UQ��8���;��~��/��O�|�����֏
�Nb��-g���,����]�K��J�R�{��m�v�E�:G54N��n=���2`Yc��Liر��#`��R�w������Q��\��-��'���_!��C�ʶ��c������G��I(xYx�,�/ӅI�����Ȯt�_n;�>j�3X�3����m��3���PZ�&���s�f��ud�FP��h���P<�V�{y�∸͋��d�"����>��m���j0m���v����Z[Y瞩oU�
��9���McV�T��������&���Y#��t�D�+�����wd> p���ؑ#��wuR�Zj�N��kw~���78?����X�(��B�P�*N]c���囖1���MQ�@�	����!a�	{m�hK<+��+^���6$Qپf{_��r��}yz<�t�^H`�_(�
չ]�[�_`��l��b�����g�� )?̋�`Ϛ�Oa̳G_�k���d��5�΅���$���G�E��⅐�Ywj��H(/H<�,��X�����#KW�]bW�͒2q�Ib��cf�1�F�y�_m�O+���4���#��d9z�����׎�gC�O�4����4�6[��D�J\t8����9�S�Ӊ{MYƞ��w���]Im��2�.��ɤ���w��R��<����$q���e�P,�CU,�>����cS��S.x�'����E��=w��i��Nk6|��?�7J��`<�R�  S�F}��^�֊�4��ll��S��<��.����]������ߋ4��^� �$�Ѡb�~�=.yh�G��<�S&%�p����b��"��+v�a+o��H��0)nr���;x6�,@�>�.؎���h�tƗ�o����Z������VR��B]1.���-@�>|�9 �tE])2�㟑4�ū4�i�v�ܟy��E)���1Q�
��`�N�WCy,�>�@��ퟢ���>��0�֘B������^���=�x�7�i�>�v�z 7Y��19�J|]�S;/�{$�\~K�Ԣ�.�:��f�o�Od���j׳j5�WYv$��T>2��E�qO��a�GS3�(P��M@&,�#J��@󤹻'�`�`��� ��Ff-�U�-������.6����r<�+������Oq�x����W�������_߸�U��<���';+u���7��.=fKˈ��x[A�ZVː�k�+����%4��6*���Q.�d��nM�i��F'��kk�\�߀�]OL�ȔD�H���%Āً������_D�M���ܦ:��\�ʗ�o^�C�tj����Nꚜ��������zϧW���H����-���ZK��*��
��vq����ԋ�#Z�e���*|���'�s~z�RL�(����"�\j�jh	l��`����	�3��F�60q&�(����2S�$�hLE��q� y�]���p@-v�?�%��y���"�x��sNn���fu��Mؕ���t��pz���؍�f� ���es\����(>���^i��H�#�PkX�҄x.�;�u�6�%�apKUo��+/b&��lq�t�*�m�c�9ӗCK���o+Q#<���0��w�0xqF��yr���'�a0�%	Z��]ඒ8=�\`!�ޮ�KG��A;�Potħ��*�2
^����&Wװ��e'ѐ�)�J՗��LP�yauύ�φ=��ht�4k��'R����?~�ћF�'E����~󐼏q�xj�#�:�%�Ց-�y��Q��@&. ���Y�2���G�Ƣ��D ���:;�:'˭�%�/�h��4�PVVĴ��,M8c�%�e���yG�1����K0��z/���W�Tם�W+G��+���ʖ��ћQDo��D�8���?��,h��հQw:V�S~x�u��z{Z[��ce����Mm���c�]�}�$�Ff�	���"J�>�q�P�i��?��dX}��zB^RrT�೗�v8n���i�X�5{��Y~�m�?��f��Bݽx'����6��	R�ǎ���>{he����*B7ę���aԏ�ˍ檯���`�"�3�d :u�~��Y$m��X�0�1�;B��o��՘���e�S�l���y�f�p3TIʯ���@�
׫�ވ��5��	$`,��n�g���RO�?��7�̠To�\��f�o�F�"%�8 ��=x�9d~%�ܜiiľ�g(h��FFF��������m���lQj��O?���\���Y]�p�h���ֽ��&3Q�WNz�T4_��æ8�n6q3k�����cc�B��K�o�-#?̐�>�ȱ�t�A�X��gE���bޙXWy�X���*_3�!y$�0Qr�%:�;�@�zj�Z����ص�Ya����q��Z�A�Ƃ\��g��	&��O8�ʲ�	/X�ݞ|Mٮ����VS���:` �cܿK�y�L���?:}=g�̈́o���(*��$.N^������}�}yţ����X8x�P�7���#e+��** {%��� H~w���Y@.�����'t�W7��!��m�>�w9h�'�[l��tYs�!Y���%A��M�x�?�ٹ�m��}��M�>��.�ĩ��D����u�5��{e��0Q��$6�b�A�H;jߥq,u�����~1�JK�dMpGJ�\�u���Սi�E�`��h�y�M|���ć}��g
�sԴ�0�y��֣/<�<�Z#'����T���m=�:�yvǓ�o�f�s�l5�wR�Χ��2Ҕ��]ϖ�N��/t�ؤ�47ޭ�n��{���.����O��~%�H�y���9� .���9��`���AE�cB?��:�Lo�h����?Sq#�<�K#��>(%Zغ��g/�UCni6��'�?���'p�}�9�h��I@m3�
/_����-֗�z�������%���e�S�f��T��=���`ݔ\�h�1`���@z^6������,�1�G뭈$���w�y�D��	�\i�4�q���6a6���33'��4;��mLR��Z|�A��û���ᎄG�e=�����W�����[*d��h+ �as +icu
Nx�]��NXP-W��ޠ«�}������pvy�|u��/��!�o��ji���8�}V�`��K=��CZC�̪r;gב�I1��n�h���n~���\-}H�偊*X%�~���8���:��΄�oh����"q�qߍ�;qZވ< �ͺQ�RF����������U��V�>q�P�\�a}��!1������<*��:�O�l�8�̓��.̶3�Q��1�
τ�ڿ���rKU��F���q����lE��� ��|X&��$��.̏����`��>G	c�N+����-%�ӳu���C��?��խÞ}���몯����3G�^Q@G>k�P���	��Rt����7���n��WGmyO�q�����p���������E�<�b�Q�#�@�K"�m����)���a�<���X�g[���V��=ZU�Ƌ3rz���DR����Z�WC�
4J*��'\�y>�S���t#��n2��$s�;�s�����t��I����;)G�ֆoT@����h��(ޯ��,%HJw�"]K��tIH�
�ұH7"K7� �
��ҭ�Jw�����S癝��{�=��cPW}k༏C��'`]����t�܆�fQ
0�(�p��.��ž3�g-��}/��u���^�h�1���)��|�G��<B�w�z )��l���*N�H�d��Ţ�D�+���r۟Es�����;�o~����R�P�v�Õ�Zݵ�@����z�eX��M�9	|���X�.�Pt}��A�^f�
�
�gP�U�G<,�i�n��QP��S���E�rDB.�����V���T�х����V_E�[���nn�P�����ږa�t��cUc�k���%Ѫ��	�T��� ���N�,S��9�yg���� ~2���BW���lλ��5\ƀ^I�.�Q���J��E��ظ���\\�{���cf�jJǭ�6�'� L�6����˕S�bC�90'E&��A���)��?�V�>�e7� kݲi��#�:uyQ�e�?S�=�D��A�C����]�ѴCG���{RO�\9��Kd)���ՃG����B�0\�ľ�ｨ/`�UnN|[ؚgӺ`�5R��L��T�_m���)�K�&��ȅc�
7�z@݀3{ʠ�Y1f�k�v��C�t�_�Lç���+��G��)?ek�IS�}L����R�/�W��nd��	o�֢.��X�\��Y���9�3M���j��#�\3��t��t������Ғ�j~��`��h���z���}��(/ny�^�fk�(=�ܸj��� ,l3h��˛us	��*[�JI?(���'w�	z�f��rr�����j�F��#�? �!w�:�J��D��L��e�6��͏[�v3���}��"ףYќC�Q�`��Q޵�: {⿐<|ݣ�֯��l�h�������8M��r"�r�ӛ_A��� I�V��n m<;�_��Vx<��`;�w�1}���j�h�����*LH�Z���B�N�сk�����YNi���������{"%���k��Ć���8�h�lױj�o�����YM;IS���%d��M��6��\H�&6�t���I������eL�s�=�jQ��t�Y��0<2a �Q͕�ϢY�(��g��#k@�=�:�_�4�@K�	��t��g.�����U$��tp��,�3E #�I(s<4���H�)?����f3��_���k�;c$�=��g�S�}�)79��gYl-�os_�dv�4(_���V-�r(���7c����������N���p�*�3$��$�+*��?�NA��h�wF�F�zt_��Ç���u����߈����^���p�}1N�t�GYz�ކ���[��bU?�%MG�N�H�"-H���n��9u�YgU���2Zq):��HQ���4��x�͈�.l�9�՚�����<�{߿��6��`���.֬��ˢ���\lz���:ڌ�qn�l��Y̙�`q����̻�F�	�~'#Y� ����{�x������E#��J:2Y�8���DX�^��=-�7%K�27o��Z:�}�?���U����$Y�'ϭ��4e=$��Q�������?��?���򕑱����vi��=�� ���X�i�%�J�EG����{��c͜F2)0,����A�/5����>]��G���p�֮v�N����(܃����.� �Z`g���g�t}�$]2�U�6꤬�x�*�K�&g��dr����I?��ހ_Q��U�6'���;y{��`U���k	�t����7��S���T�[]|���h 4}@��ɬ��E~��œ��^~�T��u��}�{��h������(�kLt'G��_D 7{A�������@�+U�f���h�b.��3����V�7�勴N����0�y����'�������)�^��D�K�����^�@N�?���O����F�:ZvC�~��V[n��>,ЬY�*/ ��831b�/�7y[����k�M��ܒ�>e?Y-A��v�'��������)U�>�`Ӏv{����C

��E íj�dgL5l.��Z�M-w��D���%�����%Λm6����v?Z��	�k�7�va]/�6<[B ����a��c�d�R�N�0����/����������'���m��R��<<��h��%�)���G��#P��c�J���^��SL)��������$t�EԿ;UE��4�L����Wݯ��s�x��(+v=so�Y0<���\qh���144��1�t,=���x�A�<�2 2����\_t�AP7���I��S������l����3{��yD7��z��x�#��g�R=�'h��+�������j����W6\�JX�d�aN��邸J��+[D�35-הy	���(����~�d��h��ϛ��`�r1_�P~�r�5���((;��\��U�[�)�?{�7�<b�ӟ�n��B��I�A`�Y�ߊc��u��<bU��	���3�UK�����ş��s�`�O������;R��� ��W���+�?6��w��[IgF���<���p�HD�*�f���v�1���^��В$g�^��!_�
㣮sib��G%*�@#q�]�,@�q8�."YJz�Y9YM�Q����>�kp'��^�3�H����ܟ[� ��$��֥�|'���m��F�/��$9�L�Q�"p,��E���}O#�:�mj��Wq(�O��c	�
f���a�X�X�*\��a�����3���D���@0>\1+�H�V7+��N�0��:\��$�t��ϦՓ� ����~.:֚H��k�<����Q���dp1�S9=b;�sg{��q�.����a}����J�L�Y5�����p���WҮ��$�aЩ���7w�8��!�;>��M��G�*�>�� �;7y?~�2�se�j�%2W�ѓ��Vpɶ c�f2U'��47ܘ�h���o�n*�2�r�fm(���/�K)�W���_�b~�����*��m�o���P��xۤjcN^�Y ��FsF_d��T-+A�ֿ�j��tm ��ɹ!i�R��Z���3�IL���L��}�2"�>�t�Ta�D�	�l��H��Y6��ق=ؿy2Î��Ex{dU�q���*�N��Q�+f>k�/c+�Is#�ߘ��(D�#>��5��9���h��f%b�x�5� � �ˀ� �0G�a�g�L�؟U�8�=3�,�q�[�2?�T���6�z&��Iz���O�\>Ҵ���}W1f�H:<���w/"a2{;"?ERl���s�	��P�jT� k@�P��k�7k���#���RY���1]J"Jsez�m�p�����߇|v�3f�ALMgի|�&�N����:Z��]��"�B�g�{�*<���a��Ȥ��_�w�H5��ML����A ��X�&�5�Kp+�D���ڵ#&I+lxK�3M&ڟ�#չh0�h�\��X����T�{�R�7�M�iS� 1n����9jj��>����̿a�Q���{��?Y����`N��'ɋ�c9KZ]�L8�a�.89���}�k9��ɇ����)E�L�k{�~R��PĶh.(�3f�|<��D�q��u��L�p�PϦ����bP�xR��2��z�o���w�1�֋�@���	����]v����i����<����W�	&Ɓ���ã�加	�#��k�.ђ �uB�x��ۆ��j@��M5ٳ8ߌ<���2�!�?��'��P�8\��'e�e�^-�}����=S��\I�CH��hAlN��tL�]jG��Oހ�}.�0���!d�]��\��-��r10�Ӱq}�}���_04qu��aBG���׏����+�*<eJ/�U�L���in�=�͏�������6�;J��J{����~�HE��Nz���i0�����Gяˋc��>�r���B�v
��S�8~�gVxC��w��I�FV�{�V�̍��L�O�/��/Ue%w|~�:y��NRqJCy7��Y��+�>_3�0�\A��M ;������"q�� U��O��(Gv�M.苞"q��P���H���T�Ӌ������s��*ZG�7�Q�n]��>"�����k�������J�Q;��zd��ؘ��I�[iU\J �v�1�]~l�*�S�)J9�����ʣ�?Os@#����]��U3<�S�#�.׶�G�~�v[� 5O>E�81�q���� Y1���1�#�~!߭��������mL���l��h�0�gg�ǚINIŃu�;b��^͢f�FA�>Ώ�N�|�P���zw�0��6��;ޡ���ˣBJc�<օ�F'-c���g<XF�~����Ϲ9;\;�C�]_��y}�Gu�;�{��"��Jd�P{��w&�}E�h�^y}]��#C�e�V�&��ƾ5���;���x	�(.�=�p�(0o�o=�u��� ����6�5=!����E�[*5[�Y ��A��9�?�w��.dF�|OsW1�:^6y�wYV�Fu��1J|��٫x�K�H>	X]xSH����o<��.@};��D�E\���$���"-��G��g����Îꎢ�\_S�shs<�Nl06%��oU@��t��0>��2�����e�.����vfuz7�)6������N6RN�~��˫g+҂�7�E*�����^���C��?U��C�&-��;A<����]�^�, �ϧ
���ܜ�C�[�&�4��_g���1�N)��o�����8��<�&����y�_5sMށ� �!3����[�].���	�x��&f�n������'G�6(M6��[��K/����a��-�tfޫ
���A��5���	��ݿ�
���4E:��X'Sdb��������^Z&�S�u���F�������-��:M�ݛd.�g��]���)K�nǦE�ۢ�3�o ��gR/uV�i|�N���6@;��FD��R�[��Vy�5��UV��tNFTQt(a��p�.ӡ���K��s�
g�B����_��ݟ�M�5fxj�t�[��BHS���N�v|\a|�8<%s�i?�ǰ���N�wS�0���Do��jFe�5'ݴ����;�����<FMo��,,��Oo��g[h���,+~��o9����wQ��-A�!�":�&��p�ݯE2��=�>
������5@��k�]GZl��S<$�_�3m�jV�0���/�'��?�,ʳ:6�H���v�ZAґ���j/D�-�����b�,fu�jE�J<�nO��گ�6����N���`��4M�U&���<��ت1��{b9&V9�8LǴ�
f5֗�*��_#�ݛs���3���A��0R4Z@�b}�p.�v`��0V���1��%��T ��`�!(�NrΆd�ݰ��	�pm���Ɛ�oJD���-	g�����5�:Q��^F�p�����o!I�ie��J�b%�������x�'�="ף��w��*S_�s�Ӓ�&��rs�h.�ௌ����H`�;�2wgӘ��gB>���#Xj�t����?� 
�y%]qN���ܖ[�*��b����O�~����z���f0j9���{⿣P����-�`���:����u�1�v�,3�7�*�;�.�W���TsL<	ޒ$cJ{�URn�9XH��=x;��	U{AX�7 V�Eb��\8.,.j��j9�'A{��_e�y����ˌ��K����K�=IT����G/u�� Xrg�0m��2b@ ��ֻ���}���SMe~bO�����;�wn�"�C�f"�#���q��[y����s���B�}$�a"m~e5/.��A�����8���c5h��A��P*��G؜=P��=�g4{����{^~���o����u-���Д�V7��|�`��/�{�2a��2��
�	g;ۦ����2�妰$��R�����vet��U�Ģo�@�uL6����\���ޟ��YDS�-ߕy~ = �����\�'�z�Z�X4U���t��ۘ��<�ͤY�uLE���8���*ޥu^�9�?9��o~;L�j��Ґ�-�H 2�L�K�J�����/鮏��y�~�[�fWVInFi�0c���萾�Q�D-�0|�y9��?
З�>��?(�oj�՟`q�]y�s�U�o6� x��6�Pf0:M��m���C���#���kS���̼�5U�&��?��ۭ
��}] �b����U�t+el��V�N(��QR@��Hd]T�z�e{��G�Ed�/�F_䤁��n�Lgݷ�I�`]���[o7�^/n�>-}Ʉ���j���w$z�U|Oj�"���i`-(����,g�R�ijo`���6̢,���Z�J�L�:�kO��5��P�M�- ��.'Y�����-�lk�	�O�Z`����vh^ܝ�L�iڕ/9h�(ۿ�D��(hKI���M��o�YV������F��l�w�������)�J��1Џ�r�C�Y���g�S�T��A��tE����S� '����&��(�tВ���~vI���=e+Gg&8mI^	<:�f)1�1G�k�AT����Q�7쳷��>63?��๐X�w��ׯ������'�[�kNg��>''A�Li@��]_v����?^h���۷}~np�w;A��_ ���ۘ?��,_��7�p��5�����e)��C�e!r�zP�`�h|�%kx�cJ����f�p�4qu�"&�
��
�Z�Ӽ)��=��_U�����}�w�#����/=@���{\�)��o���g�c�#vu�Ώ�U�f�A�rG�@+�F�c�R&�N:�4"�澸�đ)Mb���1'ZN''NDH-b:�1�w�����<��K�m�˷����(.F��1��/3)��p%�E'�S��{Pf� j�3v/I��!2�Ns7Ƅ�/kԌ���ŵ�T"��������l�,"@#+׃c)g��%cJ[!���<N��q�z}bh�|��ٚݴwf:;�1�Pa	���/�2w�V��(�:5i��� /�R&Iok ���hnm��T������ˊ���z7x2����}^��V�fv�ߣ�P�Ð~$��/q���K!��l�:B�<�'��>�ln�a�S#��pdљ#NO�l��?���z[�퍵�"M8�vQ{�Hh�������<6�5���.���FOY�����Ǝ���������J��+��w��vV9
6R�?���2^��T�6Ń0�ѽ�TVAO����~-2��$D�F������Lߣ�S�Ϛ��/��R�۠�WƩ{�H�%�'?}��ww� ~E�4��|$��J�YN��N�������C�?;����D�w﬏�ՕcT<:�`�ֺࣝk�tnY�M�[�f?D�J�b��n�v'� �$��?捕Ф�'�	����.(:�i b��9U��^�-\L�(��gzK!�����,�luD ʳ����.��;�0m����5:��}�Y&����V��ET8���J�	���R�-I������]e�;�6Gv���D���8�P�ns��
p'y��ߠT�7գ�b]�+̌�g��0�1�/����ɠ<ۂa�d�(��w�DG���k���*tk�	���Ώ �4���1�c�aj��ֿ�+E��v�$9fɝ��n��fF���������	bù6E��>��a��ֹ��Ԭ���";��<�ӳ�crd,�����ӟ�����1��3Q� OE��_�|h$�%[PF�E�	Ֆ��;�P}v7=� i�=�C?�G-�����Н�?{�Fh��qJ!eT�u����Y㱗ŐT Y��zP1ρ�ƾ'sT8�_�%ߣ�-��@����rS����x��mHI�H��(~���s�M*n��������x7��I��;��f(����E��*:���y�F!��R����d�������׬W��E��l�3ײ�q�����|e�(�^�O��RA�V�g3�oc�?C�\H�&�ZT@?t�
�U��1���5��ãI��zU��`��a�룬	�E����m��+G����9r#��L�vj1ű�y@���ZE���}��=|�DX���G�T>�D���Q��a8�����}���K��A��Ҟ��Kmp	�Ĥ���6�uY��`[9|fed�gDV��K���B$Z��uM}�AX��!���27�է�hN����*TGq�ޒ;o\-��-������H<����e�ڕC�AC��Ȃ{o}y�m�9�x���8q$�T�6��-���Bs5����N����0�hu	q7������c�6{��=m��O���οN����д^���Q�+g��K���C�~�)-���o�ǽ/������+_�3�����p�n�`�'</sp���S��]�v��yZc��d)3���,.��)~4e}}1�t�Y\΂�J<j8�H)�
��J���������;��9=ӓ	]�@���� 	 ���}4�}}����#ț#K�.��5�3͗.0A� �4������S�'���{���]���;D�U�@��2�h��w��#�	�z���Aa�Y[�*Y��6�A��3R�J��-M<<�d^F�i�O��Z�*D��3gz�R��R��u )�|�>%����|=�E@���\�K.iWװ���r]���lX���T�1^�����UL�s7�f7c�r��s��dHg�1�㻪�!��B�몷e�9���!�f��.�����O.��"��rb�?��5I���v�M7�	�w<�m����m%�Y��PA8�;���kI�-.%�h�7�{MA��`�U����ߜ��:������nql�t����E��<S��5ΰ1.�^�"Y�X�:�����<+��L��gj�BA�Cڕ�塳A�U�z��U˗�ɢ�Z��uq�C������d҃ʛ��J���5�,8.Պ;A����JP��Cj�
�^lS #2A���C�$���VkvNS1˞���O9:��&����_��$GRXd�eힽ����_v�6*��[h��#)�(���h6��^����0߸}ؗ[������Vm���'tB���ۑ����H�sz)A*�"�P������UФ��WD�R�X26�|B|�� /e��7��J�a�Y�����o9�CĮ�a���)Y}y�{S���ܐ�]x��Y`��C`����ک���=>"�JC�|����,:~�oO��hT�_�l���i��z������:
a�C���nXm���TH�½;vaB�W�Zqm���I	�ZK�y�&��H�Q�zY�G։���0)��l����W���Y.��^4���%�A?l&����Ԇ�rv���ˎ����.حiE-���W�.G}�z�Ä.ؗ30[��v݀$;��=cʫ'@!Ǔ�Q[����+�l�"��-u�(%�O��YQ�Vget7�ټ��n J\0�s
i�7 BD3a�>��N�����mɢ14�z�F��0Z�90<Q��Rڶ��V�Z�w/�f���� p�Ux)���2��:d����Q6�auY��'�(iP�n�ҽV�;�A�v����?􍖎���,\�erx$����,G���ޠ�TN �{@�D��$�+0��v�e�>CKw�2�����M��Ύ\�A`��T�{2�X��8��-R��p6�t�#?Ai�A�!���k|" `��ך�m�/AI�/k\nEv������@R5�R�q].b#�n�Nx���M� �������2e��7�/������ X�������A�շ/=s��N6���e҇d�E�ؓ��e@�LiϺS_�0n���ހ�u .=or�`&s��O��ӵ�W�pj�8�~qI�_�(h-5{&����	�ӯ�B����V��"ⷚ %3��6��j�m�kD��S&��,l�s��8S;��O�>%T�)���K3�_�Y���Yl;��:c �v���mS":~�LP��xH#BW��o�Z&i
_w�5J��/��S�O�d��=V�)=�NY3Wt�F36��y����	ؿ._��O(^N��NNv�GV������n�h�G������y9S)<�$SeT��B<)d��}��w�=�1y��7��7X@~��&�����f���.�-�Z�A���o��:*�&v�I���.O��9�
�Y�� �X_���~B�䌾��+�
�z'��P�)
j��i��p�?�\�u�[*�t��c�C������bpb8����U�R쾚p�g�m���lO�V�=q��u-��^Q�5�C3�Rxm7a������ɕ� n+�1��[Pޘ���EK(��8uq��'��V &��Q=�}&3��A�B!�ɸg��aE2:�/���@4���4d�	-��,�4�:
������1uTw��(���q��?���n��XO����h��'�%��˰��L>x���MYTϼrxs��%�V�9�(g��)�r1�T�v�������FT�GO�S�m@�2�����;/�!%���i��w���b|�fZ?sҋl��iRd�]W��lՋ��&�X�FQ%��Vrp۪W���
��^���%�.�����!�'\�,*���m{S������(��
�}�����9��wO�u����T�G���Y���,��VCf���)NW���W4��( V��g4L���i���(��3��u�s5UR�
����<�"n��B�]ީ�V5���S�'r��oc�|z�T��MW�$�hCDuìYH<	��A�r3Z��f4 �%���@XP)�-/"4W��ց�U�	�x-��׋�"#�V:0��hs��.3���Ꝣ���h�h��C����L��)�M@�~@-���2'�C��>Mu��R�F��@6�:�C2�d����l��H]�dY��N�Ž���m��m�����ߓ�߇:Iy�Y��o��A"lN�?HF#�N����;X-��^���U6��^��M;9?d���s��jL�bR�_�cxbR9ߛ��7*��/f�x�х�'�P�.ᤤl���|�]뼟ҳP�B?6�-�&�.V� �v]��wt51�����.̍�T���7���M�g����?�T����>X�ِx"	'�⪧tE9��ah����� g��Rے�e��Y<��*�5OYY=)�
�F��}�gN���>��G=�5���Ќ��9�T�0&(VWk
�e,xuS�)Q#e �)]Zl�a1�n$Ӭ���L�������5A�YO��ֲ�nYs���m������5�|搄����}k��lK���~J�B�-�l��i෉�鿬D�a }��KOz�#=`�P��\��cB=w#}�O�*�R���D���eh���(��_-�Ů%~0�_��n�x���ޑזcYǭ*j��m1g��V��e~'E�a��N�/�@5U��Ipr	��V/�N��@�������e�%�
Pw�*�x�\�'�����44�j��)�pm�3�zlܜ�X�~�5q��Q����N��̙� J#,��e38!`�L��
�·�%2a�G#f�%�Rc��u��#Y�cbV.��;2�Ͱ}�R`�O�	��p�Rm�R���Y.�J�Ov�e�4N��/Ǿ��Ԫ���l��P)#lq�Y�=k���<Y۴I�o���s_�Ǯ5�T��UFy@w,i��M��6����U�;� ��&�y2�g�!�5^w� ��)@0�Z��Y�h�T�ɽ���\1� XXUVz��I�hl����W�pU���]&�'��6����F�T4�:II8�<����&쁜��\�S !�'�Ki��$:Fe@�<:V����&	��> J��b70��Q�ņ�,��R�$��B�.KY<CJ�dg�߱�3��C��-Y����ҋ�e�2�l�O�1�t�������bqy]0UOɘ�Q�Y�z?��B��������������7D=�� ��/����O)σ;��������'��%���Y��6z��4��w�|Ҽ�S-�����8�2	��9��8n�9�k��7o�{��������Y����y,I7G')��LA��ԁ55����9�W�1J,����=�!��>�����L���Pc���`�:�=����������۟�lK�?r]�-���{%l���]x��r���'we�6!a����#|�ͷ�7/6i	�N�;�����Q㼞u=[�ȑ�`�.<�>�RPv�9�XÇ+rD��Ηa������`U?2�,��´��Gm?9-u�p(3gW��}���^�zI!)���\8{q}�YZ�;����Pۖ2�,�^����a=�M����F�K?ACV�:�{�N`�Fup�G��ū�G@�?�J�,Ɇ�G��]?g6�\���`;C�TA� �9�O�U)+`^��f��t���:��::uNal�Ї�D�
�	Y���]��IG	/�+`�:�5ȥ��͉$�w۸x?pE3�J���n��m&�B��٥��B���S	ȵ�/����"�m<?�=�x�a�܆p�4�'A]BH�8LR�>�MQ�픂I�`����<puU.�����xYAӿW\ � 8o���djڐ��x�z�Rn:
fpL�rYy:�E 8�_��5�C±�~S�%x��Y=�A
���	c����s��#XS�N>E'OD�b���h�u��+���bc�G�d�e���RRK��(5�[�����<��An'r�c`�E�9�vn7�}B<�Ш�[U��s����'V��o�4FF35�5�W����UPA�A�-X��w�et3��3hA�g�j90*���#|M� ۊS��ѿEN�5�(vE�țJ��{��W�g��^(Ď&ۓ�bww*!�M���`�.�N�����!C���hk���fL�)Z*_m�B�-�[G_���R'C��� 7�k��k"$f%�f��i4('��Q��^�m��]�G�"�	�l|�M�#���7�y!A�:� 䗃�O�������f%_��3Rp�8�]�S�0{��V��H����Zo�o�4L�>�GSJ�[�&��Ps�0P����yoy) ��j}OǓ�BB���FV��9X�#`��N;�����E�\f����l���d CZ��|�{v����6OMė��(k��y[m@��Mi>��K��0�Ƒ9����0N���2�����Gy�u��;?�-�swd	���~Ķ�|��iE�?��T�����QW�;��d������Js���Z:
G�f��R����>�j���"S��Zn'��`3#�D<LJҩ,�/��We��[�
"	�P��M	��_'��fRS#
�:�;��+sW�l���M<��w��iOq��G ���7��E=˻�v�=���L�m���b!�$�'�o)���q#�f6i-�{t�,�� vCT�n�56pV��pb����4���5��(B_��j�a��8y��}��
kNU�G��G���z����O>q���������$��B�w$���Փ��N �Kr��c�������Pa,���{���x�Y)�]Ap[���c��?v󁞆����n?e��B EM�}�i�'$*�#��X��k-K�k�ڷ)!e�d�b���CN��s5�bn�l̓k�������sϤ(��G�|��34��/3Ƨ:s�+\��kS�����,WD�������e ���G$��< ����V	�}5�t<f:������4������,�s���4����c�g�Y+..S�6Ak�&�L������幪�+J�y�ƛ�2��'yx����|*~nɆ ���5��Vw�R�:$�< {I K��K�ܛ�|����|L��r��6ާ�o�2>G^a������1q����j¸~�����۸|�k4k�󅤢�G���J�){єA����^IW���w�n�cuM7'�Q��Grwn�r��S��������w|N���ڢ%��uM���y+�ί�-oW�i����p�8�m��p�M(��Z�*��(5C�H�"I�c��0?b��,La�AV��a��n�D���G��(O�wqYX!D�Y��g���7�l�0��	����.��	k ��p}X��C���1����t��O�wj��ͅ�{���kB��n�w2YѴ�\l�	b�W��y�)��x2a"����GJ�*����`��ay��%?=���e�lZ�{�]&�����Y�@����Ф�]��׹�<op����Hp)3�I����T�l��������|�PA��m�0)�y"r�e�s ��ƝW��S���z�~J��Ћ����Nݍ�$�C޿���+��oKX�:���w8i�ߨNX:/;�E@%�{?���ڒa,����6+�V@$����&jW aub���@CM@�|� �����/�р{6�3�����Sn���<Q����k̄���cw�A�x4 ����rVgR9O<2��m7$�p|ґ-����bț�>[
�.�ƷM=o���@p��4���'���9YH4��ϯ٧�?�?�(=�4�Xb�WC)��ռ���-Ț�L�q@ �|�5��_�BT�).�?{�[K�H�
�ԕhB<�:�n���# �a�|~�$�SP�v�-+�J�&��g���L��E�ob?���]a���t6X�7I^�m�?���!v���	"�qDջ�B�nb5.��$�ג{��i����e
MӜ�n\��GS�b^~��i�͘�����L���{U�aQe��f�,G[�3�J�u�K��2��-s �_�K��G�ɞ�M読��,�r�E$>~��y��h���ӏ�9��s�bǗ�N�!��2{j't*9w/G%�~������6>1-��D���ΣFA\"s(m�1*�6�3+��x�X�^�"{��~ �����KPc�z{�,��B��A�	����$a�/;Ȼ�J�JT ��[Utsm*�U�T?JY8�:�����g����K����1㾚RW�=>�Ds�F�w܂OL7RA���f�;$��(EE#3���r}�DR�g��'���
�c�G��t<o"8�D��� �����3&Ff_�&��F�zJ��mV�WK;�_����td�L��q��Ȇ�MF�=q:�z�B��2=��JK�R A�������v�V�ś�׮�'�����9�-XJ�a}%��.v1:��	c}����`�y1ä#�ݖw�q�ڎ�ǻ���	�G�:�<�����2�c��m��G��6��e��LM4e��?E��x��V0��j�^f�����GMt���r��|�+�8zʁ�w����.:�	%k%��ց����Ϩ�����?�i��@+�f��_a��Xu�x�?%�a�y��tF!�l�E�M�����n����s��'(��~��ƋG��@���A��6�TL�0�4x��W��nrq�a@㋗)-�8�s�B�r��1��j�^e�
��2�y�ɫ����]]x�/3�	,����A�\�G��g~[��`W#q��2BQ7c�Ef)Q5�}�|��M���]�����kJ��r\��	��#҃|ֈ�u�7�sE��n��#��2�J�8e$��a�a���Q�]����a���@�_G�	U>��y��Qðr��0�gq��^+K�O����D�w	s@�
��Enz=K w�[dk��7Y꫽
�t��V�47@DL�q�ҹX�朲��;$0���e�Ł9�����NP�іz̏��`A����Ư�!X���%n^-�����9�8��S�j�\�6��W@��o�L�P}�!�B
�����]��ѱ�ǐM��;֟�{�V}��/xI��k��\_`�/��I�u����C 'f��L����y*R\�7��H�����d�x��ǭG�����룢�	���7�-%PqC����jq����i�%�Z *���b�w����/�-T��قM�y,��l�տ�x��6���<�P��R�%�~~�B-�	���?�:j�����\)ȶ�x�q�RsW_�����׬V�'�[n�H�c�]V�ͳ��Q������X����7��HQ�p���;߮)�q����Ƈ�������e�!ө~�B��������[j蹊�����ٞ�>��ik�5�l<��sV뷿�������vv^~�����5Efy����lt�@���Bqʋ:m�Ao++���yסy�_����
�&��2�n��z��u����ˠl<���Ro(�l��|�R�����
f���#�в�����̣}�*������}��	;���sz�t��Dc��6"Ž3�y�i��nKq#Rx@B}��k���}�h�u�6t�Uj	FL%��b'�O�;`#�ۋ�ΖR$bn�)>��9����k�<�����ZX$�F�Y��LN.�|v;.���b>����!([cf�ԏq0^H>%{�`,��c�#�Pn�D�wl�kn��6���ȤF�1�i����_�o�v�H�<<������	��C�<�7=�wd�A���r����ǕI���������V�ϧ�J�+>�,7�1��-zgQKGGku�Q��]��k�2� �B&D�V����b"��q.�Ǝ�����;�f]�5�����Y��e�����̬���j�)1^�%#�e��������=�|���J.L��m��P}Gj���$���;`cﱂ$����u�bSP��f�V~���К�z�E2���1{���U}	4���?�H��[F�H�De�%k"�Ld�$$��H�]D�.�}_�$d	a,��2C���G�����s������s���z^��=�(+)��)��w����U����s[��jӶ�Z���Eu)�@�ߖa֒?p���Ν�ŝX�vr�y	8����+fn�w������?)�O�J����Ka]ɸ��Y�D��z�R-Vc�k�|�&�zDT�V��c"/8F�(�5Mdg��? �/�Vy��\���233{�Q#]%i�����+�l�p�3v���ſ�D^�����HU�I�ܒ�A���W�L�/�����������@.���[���.�o��t%���t��^��� ����u�~������j�O��� ��&BҖm�B�����5�\�ث�//����fmwU���p��]�w�*�$H+�(��m&Z�x9�I.O�z����� ����rejjW�c�l��et�S��u�?�7lKc��|��j������X�.{ْ>�ҭ��w#&�/�Gw��Qfk	^��xa�YK��n�]K����{[�V�}Y�JNѾ������/�o#�W#�����f�qao��\��Sz�}�?��v>�Y;����Z���)V��L�W��.&EM����_�;������xNMl�����4z��˄z!�D�������R�r#)+g�4�M����g
������_Jm=�)��f;q�{��UOK�ζ[f⎳�>��ؽ)!�#������F�銟�Xf����vU}poP|SG�7��Jm�=��%	@�c	�FC]��n�^��j��+g˨¤$���d޻�(Ч�{?�j����,����G�{}e����Kl��F9g�k��9�)��ǵ7�E�(o,_���_�� sow��O�s�@~� 2���n���_p�g��_��Fgk��h�5r�?v�.�d�n�E)Zhx�������:��r\Â�-���j\�}�?RgӐ؏=[T��8���Y��<E���_���w@�4�7Ƥ�O�,�>Z�����2����l�r�r�D?ػ����L�F�Md�憧6wvv9��fݩ�يz��;6Q��iu"`!@�oaQD�]Έ�~p��a=t�i3�+V�Ŀ���8\^� �;����^U��G��ky!$A�M��L�i%�N�qd_v�aJ]�LOeF�կ�s����9��Ú�Zs�����c�>eTԕ����/yC�c���;|��z��cɵ׫�W�Br������<�������E�
s�z���[�Ζ�^%�5yd�a_t���|x�Y�鑁�ʑ�-���_"�!-	�!\էaO�l]TA1+�U>�Z�;�L��)�_A,�VZ�������+�F׌�kn;�-?w�
�zQ��S�=t��D����#/X�Y�_݁�FB�^��K~}{Ah��"v\�D�n?7���b)�b��ӊ��E��^����Ʀ�V߫���:/ǰ|s�	�h�i���I<Y!|��z ��[T�ޢE~���zę4��K���R�|�Ye;^���d5}v7�c2E�$���/��N���W�$��+�%���6���d�2��5���Y��N��~:ĉ.��BU�{������S,eXY ���"ֆG�U����3��χ��� v@f�OS=ܛSn��\��⵶���Ȟ
U�U���ۋ�����\��UQ�#��>~�_�+��i����ab�{������Vz517����O��O���VKi��w����
�&Gq{X��J���`U��zq��+�e�q��h���
�<|q�^��՚��{*;��y�����ό�Cn��1 ˀ���sג���(�?�(�|�[��~u+O�):����(����-��������c�cu%�ҵ&��u�x&��za�kzw[����̻�<�
-����YQ�oz?D��}&�Pwz��{<m3��h9�������L�.��/�$��^Kh��q�Z�����Rm�ңb����""�kWm��(��D��/Ge�Qx�ӅN_��q���Ω��U����ߝ=-�Eע�UG����ҭ�If�Ԃ+	�kߴ=����͚�ҙ�8`d�����FD��-.�J=dz.�\@�.�T���d3�
��g,~��7�%���Bb����[Cs�Y�v�k��)C��(���sLo|?Qu��r�6@�e�\:0�3�i*�>^��K�c�_�{ƳZj��HQ~�{�=��Ј.�� ��|���;'C�~�gq���1���VTYyA��E��L���v�����ttYfc�DL �?��VU��5m^gTż��˭[y�������*�n��	E�}���F����F���*�vɞ���۝�
P��<�ܛ�s��;oF�Z��6>������*�04����}E�cZ�=��SF���b�*���x�N��׉ X���6E�mm&*iHk�=����a�X�=��`�~�I�^�����5;{ڜ���J��fR=M�]�T���~����v��k���I
j�y�B�=4���e��>��Ii�V�)Fٟ�+��=��a����Ez�O��Ʊ��!���Զ38kc�R�G'��3���Ykm���?�?X����5V�(����pJ�O��]�aMb��8�楸\�x�Ey�e�a�a��3�H�]�-�+��~5za+�3�er�/��xw��g�mVR��̰�D�����@ps���@%����%��L_Z�1p,!���J�q~�s�l �o��M;Q i�W�/x�֏��2ή��������U��P�G�ttq�~�[�,�z���sox??;��%%6�D�ύ�j�`�I'�n�
n8�#b�7����"�P��/`�ڄ�9O;:v�=}n�f��z^x)��!�s����&���!����Ղ6�f������ -�AZ*�$�(�6����K}�ک������l��[bN#�j�2)(�[�j`��,Bg�cUA-�=݄O�ȯ���f�]^�$��]-NF��=�/�b�Z�o$H����Imz�=�w_$�?"�psi�sظQ��B<��9%��������e9��)�y����/N��ć �w&_s}Zh$ꞟf
��� ����dCc���%V����+S�yv�!ko�Y�~��=�F���v}�i�`z-�F�V`�%"����c�d ��.|���X�pM�cV���\'dAֻ��A0����y����;e��4�mTūPH������	0Ɋk����d���\�~�5��k�B.=�:�UFʹ�� �!����b��,��2>EΝ����M��<`������ݹzM�;�Їp=��׭���!���WAy��Q�Wf�݊��,u���\Ѭ �Mo����x�'7�Ə\D�Ib[?�X*3��q�I�\�M�xz&d>]��N^���H������.A��I�-��ߑ�ҵ�ZY�����C�U�F�)��^�N�p�;�
G*�,c��=ѲL:��B��n:=Q���dJ��`���t����^��9���eKZ��Z�/W�2�Hs�iLk5�d�;ib��U�
�,���]8��ѓXO33��"��-"j�������-���l^��=�و��3����R�W��W�݂��-�t�bPC2=nyQ�Ց�g����I~�PmV�"
�#b	����{)s������4�I���M��@�]d{{��*���h{�|�y�Su���׾��K��t�F�s���Kym$��]⎞����T_��)T����ެ$�K���I26����O>�_�4�E�g���PP�p�? (�h�ˍUs��Z����:((�<B#��S������ �:�}p7���� 6U$�B{�@ltV'��`^*�et^��;?����z��ze�-.a��C�\>Ù��A��jt����=�������X�1$%����ƨ˗QR��n����?Q�/�������.:�|)\t�m�=O����-�̀Ѻ!� )	&��qB>V���ټ���V�{,P�}t=�d�����PL�T��M��Z�@l+��tt�M	��/��^$1��K���j�0����������Su��/�_���}��]�)M���I�����˓�%�啷�Ē_�;"��a�?K!�s�'��O�}*�x19A�fl˙�WN�!v�uw��H��PH�@|�p,"QH�b���=y#��sD~�p�b�\��x�`x�k5Z.�����j�L!��-O����B�������\N����W��Ή�MS(��f8�!ѓt�%����� �rGc��M\�/�\�7w�]��̬��gkտ�<�e0�����s�7Y�+��]2�]Y���4��k$4�B������;�=�d�-�|Nr���8�����c�d�H輎�"e��ˊ��|��bOnN��3�ogk	�������L�j�!�g^��p�g��-���a<�D��-ZV`�%�{�h�C��~`ӈu��v�\���R��{#ίt�W֊2�s.~��B/��M���^\�I���`/`�:q�O.���~{�����M�5���2�
z��Z�ū��F��oQ��R��4�<R4�Ox��HM|����L��F
~__�f�0>������,��2��� �'��?�1����>l�Y����wAvz�$i"�'}τ̌밧��;���)��F	�a�A�8�o)��緟]���gi��	s����k��A�k)��ʒ�r]�Q�k�w�ޤ��1�v��Z8M
_�3�Hw��낍xI��[5z%"U���'��uB���ɱ�,���]G���RI�0�xP��L����wo���+[᪥9��N���˞K�/���w9®�O�yX��:����x���R�>��<��j���1�őy@̔�{��.6�Ǭl�Cny�����::D,h�@~�;�d	l���W���60���Ɨ��F��r���I�?t��2��H��<Y��d��&��;~���G{��l�,�u<�˗d�#ܟ �	<V�A:9�Oi8>WQ��m�}�8����U+f2�V��g�&�D>����˲�\��9��;�T�3�ϳ�X"�n�!Q�Ldz�  OR���+�J7��50�/�S�N�DM�����Cq��cbc�z�'
j`z<�v�D��j\�G�}�*���d���: wu�?��a��7��^�?����A��	ÉK5��yWB�n��թ�Ur~�7	�AZ�)��P��&x��[	X�קg«|����L8ʞr���N��n�u�x�;��#=N��B�E���~���GN������q~��Mg���Vs���DZ�_���X�W.���IX0���텥�]��$��7�㈄����p��$�O3@TKi&�L����Ej�ronS3"�n�.�b�K��"8�����zҋ�K���D#��憏e�P���	R���"�l��;�K�G��\\�6�w闍.��NVi�l���+6��*����6��<>J�P�f�+n'�.�{�;kh�H�>��BS57�y������A��r��?[���	�X�k�C+����g�_�?�(��{<p$w0��6�2�fZK�uM��3@�KK��	��+[�OZ����]�4�}XI���N�< �"�C���4 z��	��%��Wv
AV9YZ���ʱ��|��6s����ם�8��/�լ���J ���S�⏛U�oė0�X�[����wD����E��u��J�=���++g�|h�	�Y0%� X��F�6�P̛�ę�Cm��&�?T����`)�rO�,���g�5	�����3�����m�:i<P�I�D��>*W��=�u��-��cz15�ۏgmR�	��8�С�n!����n��5�#��~0�[��P�8Nw���¿qN+_[��|2+�=KXI@�)-��h��J���F�����������=P���8F��|�����uQ�ܠH68\%�S��I R'Z���R�@�9�T��*~��0�xb�:�L?�>��a��J�5jM�RLpi��"e=T'//���?6K�Ptz�7׾�N�I��f��0�%qv_��%k`JC�-�g���X;�N[и0.Q'T��Di�"_���a۟�aR5�a#��ۥ�`�q���'ލ�I�`JU���}�h�����% 1@ų]��Ne.�J�zwV��CR�����;�m��4#�{~�o^��x1u@Ƕ:;��b�x �3}�IDa�O�f�RNL��/7+1�Qs��J4g��y5}�NTNu���5г[��V>�	է4.�g��i�S�zB��5ٱ��L8a����0�����>�X�l/m.���s�_�lҌ�,���6�M7�*��X0���Ĺ=�Ê���}Ξ���) p����qȅ��~��	��J��]�r�n��J��*ڰ�?˸��{�y�σ�?��н����+�����X��`�Ws.���#r�SfBQ��oPD�UɃJVg�X�=R��|�V�6�����
�ޓ�:��䳏>�۹s��ںR:>�ax����D�6���Q��ZNx��R���<<<�9D�4�|�0�_���-f�v���$��s�e�����{:�E�kfV�h�\e�ƙqE�~��<cUӾ��7���R~+|��LR�Z1�v�.��v�u�����;u�gീ�v?�Z%r�ґ��C�x��6(������>�)�M�}��3A���Z��4��D���fq�GW����"BFB9��@WH�� p7Jw���wz���E�o���8�d6���hj]j�X�ɕԸ���o���ՍZaX����&��(�ݠ��l���$U�J�t���cA����g�rrF�,e�&Zzo������(�t��s�:6[5Br����5A�Vu.'��6)��S(�>�;�K��x��Ã]�D�x2�	��VNa�/�%�1�9�7�%˟�d~��.|�:3��Ws�B)ۓP:�?2�`&�q7H������㖴 PD��J�m�ְ���������_��h���},��pl�-=��+����'��xf��F��=�_��ͻ[�kP�fx�i������*k��0�k�wV�^�=��sɏ:��2NDf�+�����a�q�	vle�}�.��������w6W��}���Z�PՀ7��b������g�=Ȃ���]�68v�������^I���)ȕX��H8>�w:��<��(��1�31e�!_�e\w��4?�o�(Yc�Ӱ�I�����T͜�ݕ"���� ���͚[� 95@������5]z�kK��b�6�s��XT���$OV�=��Sֵ����_��`u�n�{�S�Krf5�M'���blX��h	A�x�(��������(��:Q���@;��I[�|5� v�`U~u�[�u�?��1�Y�M�G�p��>*�<f�om�IE	H��y�,�{3k3��>��s�܁/y+�,܂�gk��UA6�z�:��ɮ���,@f��$hu�ېL�n�	tZ[�p�|��(a}:���Y�a7�����43��(�}0�½a��T:1v�[��[p�r	���'V�.6Hݣ��k����:'^ٖ*��CvF��l�Q^��Rl)?�s_�M|*f��0�����'��H{Q�h1l� ��p��Ců��}�(|2�����#h������fL>�gR�B��mz�μl�
}���Z��@���M^m�=�0�8����>-�����ot��M��.3�A$��_(�,����ߒ ��z����4i���gӁ4����7�[]��3k`l��eA���y͌�9�$�t�o�fe�@�՚���_NT��n��{=V'QרP�n`
�]�ek��S��"p��3�]=v�t�a�1�d���O�VWc�����{M�K6"9�i�gڲ���N1�����\Pd����� ��)�_�l�hw~�	�ͼ*��鼤rß�����Ao�S��y�F]vsp����_ٰt��� �ǐ7�
��8�3�Chr�%����W����N�540#�q	�_�� u�-}g�N/���/i�f]���S�6�K0>�Q���S��1�PpC��HH�J�ר�Z1�5w�^�B��~���N!-�\P�����18+"Q��#3�{��knk��L+3��<�n������h�s���|d� ��Ņ6�
��P�6�r�Q`��\;C�u;W�r&��T����ߗBE�uD+���[U���J2=����*j�TfBj�F+<��<�W�rcSI�a?jݻ���ϒ(<̉� ��rO�"��!�}��ݖSW�jdK*���P�'�{��QC��E?�]9c>U4��L�n�q�U��1�y���W��f
�O��ۯBr+mn�,zm9�tnEX%a5��̑?WB����$
����ީ�����wj~M�誌V�=����u}���	�-M�Ʒ�W1qU�T9r�\ ���Av˗�[o�fuaN�n��5xgV���@�<d�9\m���Au���Ǭ�!N��>o�Ӭ�T�^�N�J��� >���l�=�d�V}�:n�{���x��rԂS�X�t��T��$�)���ݗ<�|�-=Acn�ֲ-�?x2��恾�Y?B-�z�y`��E&Á%��ԟ�������}�&�23��3��5O~�ǵP*
��z\�~qM�����cl�{wrn�B-�W	�@��J�+�A;��ϴ�~V2G�
ފ�ч4�u���G,=J��K����(+���e���P�B��_�vy�B�B�G�������<70�?ݟg������a���8wF�p��Ցfuj�{�sa���|vӒH�WM-�<�>�'ob�&��m�&H K��cɈ��L?�ě��dx�#SC���نe/�n9~���q��^C���×Qp�n��H�Gn�r�5�^�~v������N�iVn��MrǫiO�o��|\��Y���;�\�hp����ł�>�{"7�K���C�X��)ց��XĠ�&��I�����"�M���CDaN/�� \�����t�b�ƅ�������Kt�LʀE��=F�5& �nF����DE@� [��N^Ǖ��H��L��t�E�[����`�ΝCp�֎k�`�K����+ǫ��X� A�]E:wɓ������C���c��7�&���4��r?`&;�8M(:�}Ǩ�5����@:�	z`H�����Ok�����,X�ںQ+A�ID�$X�HT����>��G�a����d�QG�!�4�<�:=0Vn����HIM����ǟ�:�(E���X��Z:�R��t֍�����Vz�9}�%�\���rvz��4�H�\�D�����=![��șkl�n%@�[�(<��z�9"/ޟS����EOp O�#��l`�n����?��IoC�w�[�0Ab��p�k�7k�1tbHe�
)2����&�����X:�a��N87Q�ؚ�T�����Q|M��i�� P ߤ_��)yT>:pYy�cB���J�*O����*g:���/����[Lfݩ� jck��Ũ�=~���Y*���u�Ѱl��T�Ns�P��]+ǵ��^(ZB!')	-[�s\�����0��Kw�R�Uf����`�%O>���Q��~X_�b���+��g3�ʙ"RZ���W�\�,��k�x���3�u0�5E&;_@s�gGTl�o���=k�JB�)���Q#��%��h�qz%�f-����n	/#��@�pX��'�ou pW�;��(�l���i��K ���g��������������#����k�A���Le���i>��&'"9 4���v����; ȕ �]��P�f,��	�5Q���/���D�/��@=��H�X ��r���\����\v$r`�֍+�C*25��`�xa�R�f���J��ŷ��LD�]`{h�|/7���ֶ����p�M�.t����2O l��1�/�|�O�j����I�ˌ52�ˇ!�{�Z!L`���&Z4KLȻB5a�禆�z�˗�PK   �M�Zr�>�� � /   images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.png�gTSk������H�o)қ�4K�
* UB0��A�J(�E�RUB'�P�I�ރ&�jh!��Z�����1��{~|�Xo����|IB訝?�v�����}�m%g̟��'�_~���p����O����s������\�����Mv�􁇬n����m���\���p������ճ��b�.��k�lTTQ�Cn?�LY�rp���M֝�VOY��u���h�~f�����y��$+e�%+��2I)��ywK�*����ƋAg�?��+t^.7�.p&��NG��wg���~I$�_��i�"�pw�e��͈�t���47w��x�[��� K��ӓ6������Pu��ʏ�/���Aa訨,��x��
3�Q�A�4�ɉ�U�5F�0`}��{:p��$�]��I�ץ"��' 5�x�!�A=���=����_�L�M�Jj��*&)�~4�Y{�o������ }@b��D���!��/�+�M��u�5!�;,Fə�@7��jv.���ɛ�++=w�-Gx6�Ǎ�'���HQNS��:����>�gE�3���Q�Dha���^�-0�[��U�����/�a7�Z�|��d佉	��޷AL ������&�`HU�9���?n�}��!_d�Y�9Ҭ�	s
<�w�Ԕt�h���Ip?���T��.���ͽ�W�:h��Ճ�P��X��o�N�^��n-Nդ{�b�/4�՟��σ���zG��`�����%�&���oX%Y�*�!)��#��J&������s¢zG4���%��(}�����GY"�G2Uץ<
Y�H�Gh4��'j��J����6�7]��	�&�!ٱ���u�����Fc�4i��4=�1Z=�0�޸�/�X�X� @�F�����Z�W�q�8��ya>pO�7R+�Щ`cc�ű��8ȹ!7�ly�<)'iQid�LRc���NaUa�7�Lړ�����#N�U/dX5M� ��5poO,��w����5o=3�奚��mm�U}4),��Y_���ܳ�ߢ�"dе�F:���㴊�z�F��U�E�0t{&����D4���M ����J�;���x�ϑ���]5SJ�7���a0�Jvc15=�or�}ʅ�Zٻ,�*���}:�Ѐk�^��~:U!�1���W�Y��cuV�`�J8^�m9���@����tЛ���8q�v��7+��8�����)2UH��P��@vE�v�Л��{��}	�%0f�H�"�9? �L����{6����n�?g�\�:�1�#�{Dt�f����g�����pI�t"��۽���d�9��H1��`F�ܪ�迫���>�E_�y�5���tz^����s>5�5�q�^�0߬n�u��k}q�*��[��к���,(�7�JɌ�V^x��a��^��MW�Pt��R��l���Z��,���e�-�I��M0�.�����۫,�c&��*�C�9G�M�;��v@(g�rw�5^9���7�҉��H$RRq:�MHF��c�?���Hy�f�X{�<�!�;��g����\z�nvj�s�ժ��*%��0��+��I�������z=F#33�����Z:�#��*�x
>]�0�������C���<g��6D�1G��f]�$��>�����K}�|��v%��O��:��L�|��r
DĤnԎ��ld�Y��맑{�����ޔ�T���Z�v��
�����2�̶�ݨqFάP�ԧY�=�܄<�|')1T�!R>���{�����0�;����K�V�����<����	rq_=]�*����n���*'=�Pg ���g�~v!�y2b=퀕.?v�ui"@P4h�z�|�j�Y�u`�xvx����<��e��GLpo��n����5���V�ꢃ:�5�U�H����O�UN:�O�_���~�)&��Cؗ��&N��.��RsQ �oe�^����h'5}�k���?AC�!���a���'n��i(D��*���H��Q^^���x��qu}w�����O[�Fsz��ir��&�/%����x-q�.��D��!�,���@���= ��|ډ�f�I�׬h�)ĂUI�\K`%�*�1?=�UL}���4\ͅ �~��N�����x@ !��)���}N��z>�e7��>D��19H��md�+����8�ſ`�A�#��#��{�CY��/���!b����[wÂ{
�,�"���د˛�dQ��x�����0�*�t挃t隒o.R ��"�WQ^�6��6���u~L��4���:V�B|KP�����55�7�#�aQ�}]ԇ#�kY=��q�R�����Fh��❷j#C7kF�, U��$�_4S�������wF����ۋ���4�G�iq�:󪲊ѽ>6h{�eF��V�XA?�^�c���^��Cʁ�F�.x� ?Yc5��2�V��C_����7�`�RX���(���Qz�����d�7�)q��S�4���GARzz:��+�����#�j���몚�%Y����a�I��*�`��1\�Y�>�Q�IM�:�U"��Bkٱ���.X��bow� �������������� 2�|��=�B�ƹ��wU�k�~�����x�������_��B��H�A�r��¹��P�%
�a�S���NN���`e
�4b���AJ����eI#,�q�;��������<�(��b#�[g��v&n���j*S��	���
;��V�ubM���w��Mi�l�2YW�:�Sc	�����~�i�}�����xN��U��ѺQ�c�mV�%�4���ƪ~=���@"�I�/Q}����
M���x�2ɡp9)
��9����TĻ�:)��(�$�W��Daa��+�M�A�	ѳ �~���ď�
�"WC�3�z��G���{��@T̷�~���}��6����JPu�C�Nܛ w0�76�:�`?�Z��x;�Ta�W���"8�#��ȉ�)D�<��uO�u���c�B�u��%���XOJʖF�g,�������*%b��>��N/��������N��HM�WA�4��M�n�H�˫��U��#%��=(>��`j�S�Dd�]4\�K;����U4J/� �6�# ��x�{ͧ�ۋ�<v�����n����vuu�ۭ^�w��v�ᴗgu#t��l؛���fұ��$~�1�ytMC��p��M�ܴտAx-��{�i��8ֵ���������B䳣G����߳�(�; �!Fft� .?��Λ5Ҕx<�y;k|s���&^R$IQ���"�������zz��"h,sn.�C)�d�����H��O��X�0 N	)=�%��d�B5?w�Y6+�N�3��I��2c�q�05Ymԭ�F�!lOR������W@�X�t�Ͷ���ۥ�U�R�X�-���B�OVL���6��ᨆ�
le<K��ӳ\�����_ZZ�RϢ�F��ue���B�<��Y���'��{QB�\��&}�Z�oա�Ǽ`�Xz���P�KZ��@�/�4S�����3azn��sd��MFg*aYD�pZ�eP���}��97��t���y5J.3߬J�P1*�k����t�0�Fadg�k�z՚}1�=tӽ�5�v��<���/�0�DH\h���ù+����*u��u� �v�	��X(=�G=�x�<�U�F�2Hu�l�L�O�{A^��@�'�i;��^���9���t�&=�cK��� W����N{���,�~���J�G��!�C���E��׵Y Vw����z������ĎVY�79�'����k6�_7,f�M�"���u�<oM����$�<�.2��Ë�l�(��J�̯��@j@5�H�DO��[���sp������_ �(z�� �?����]�=;�p��un)a:ƭj��d晴��W��̃�����R�r{�\=$qa�ȿ/�~d9�%i���6����ON�",-�<�&��ڬr�mU�7Ψ9Ց��׏�I��X���ǻ�޹�KJ�K�X�5��2 d�J��!�
F��a�moDs�*Eێz�~mL�/��w׌?����ܱ��t��1����!%�As�����5l�j��f��ڬ��>��ƌN�Ƌ�n�&bJ����W�3��[7��Q��:J��\o�-�����,5ܿ�D�m�G�Hሂ�&����I��G����(��X]�C�Y��FM��ВIzzc{�j#?	�ze�u|�{���2n5�CaZ	�*���uϞ��m;u��Vf���[!j6g\ax��1f���J bwR��iF�&��f�pd	(���a���?�.��_�Ά����{f`v�Q�3��Ī?���>Y�"�;�h!����4�}/9L(�-WHs�O�b�8���]� ��u0n�-o����g��oZ�J��x[@�i�ajJZEO��0�:�b#�����dL��Uި��"m�?#�<W��`Y�����՝��}�0x*/�ͻ�2]d�Z[C�c�/�Q#����W86�]��:�N��L۸�w^����f �7iʃ5 �.���쳳>�L&�E)���O�x��̥%R��c�N)��!d�kۛ��P�?�pt ��+G���L!��c?�U�M)Z�>�K"��@[^g#���X�iM]*k]��DD�,�ظ��!��WVt\>�I#���[�2�?+���u
}
o8<�[��S��>����m'"@�g�K.�1����B����I$���RY�|�f\᭸X7�:��WFa��(���]:�� j?���~�����G��e��^"Ϥ��? ������y2z����M�ˢ�+j��Q$ٓ�ha��b(1M��Q]�I�t;$$=�NQ�~�Z�FW��� "��QS���N�Jð�l�%�*�X)~�*�q�W����ܙ�O�q�D�$-��N�5q��dk��oV�������Y� ��|���
��G��6�!im�+;;�t���*F�="$����"��̠��6����ƶ��ĥ�ɧ�t�n� ���VR|����������J�Ϲf]�X����G���C;�G%����?�;K��O?��6|dy4���r3g�;>��f�2����$J�zՒ�M�d�-d�q��.�����!�lYi��=}��{`��v��v��(�����H;J���'<556W5����{si��駕Fn���&��/'��u��5	-�F·������?�g��`�_�g-�;�	��H��U���Q ��^5ЩE�
��/.�o����'9����>d�א�vr*�}%l���I��@�zP�rD~J37��):a����@fr��e����������w������?䖿�� ����m0��J�a4L<y�)M��qc���_'2��[�5������>	�]��j�޹P�쨙�s!�_�F�W�s.�|�����?�]v�{D�x!�N��H�)�DKK{�^�&n*N���h�=���$�g�|��ύ)7�.�������{��yQ�nY�eJ�P�TP��.U�U�g�W@K�z��z_����w܋�͛?͛��̤�[��3hzr��U�L2z9�[�Ϗ���as���Aq"�`�q��>6u>u��#5�
�2X�O��>����h�*�*�W��߻�P贆݋I�C?z�fL��X�sC}Sna��to8�8+Xɽ�A��\En�ʄ0f�gG�B���U_z<aȠ��cPs3DƮ�5�h�r�}E�{�	�ꎿޓ4�U��j���=�������?rZ�a���ѭs���iV�W�����lFDN��W
H}>��\a���`��=�I	7�x`w��_��U������뵳2L������'�+�w\�٪T�e����[����W�z��;��"�VE4%FDb��?iѮ��xC*��g��z�h�]�pn0��=o���i�{��U7�TQqq|�LJ��۽�K-ǮV���ry���o��+�u��h�D{���?���7�zo�h�j��x_�_�ϵt����~Th��Z�����ͣj��="v�H��Tq��z��k漪�<�����b4��
�w����f>h��֫~5Ȍ��g[lg�0���WOnn�>u�̵�h?x��j�o��*�C7u�f�T4xc'��/5SvcĹ�Z_�%�L������A-����,_kn�_�e�O���L�^���"�{�S\bmv��h�1͹�� �~�v���3�i1�'���l��l~z����.�nM�u��J�G@��ݏMO|���H�f�+8|�^[���K,���ӡk���1���_ھ_�!`X�.�Fh6,�(dG�G"Hx�ұ�9����C���+;+��O�""L������"z`ߎ�E�`_U���^"������u̼�B�#���鿎m�u�.[�8q@}�:=���whb�N��V7?�ɣ��N?{p�������
��(t=a��m�3�/L��}��V��(�s��"}�^�ıe����՚�PU|�ޙ��1��t���0����9��ζ����Tc=!�?Y7m�g�R�>>��fڨ���6e���r�8An3��N{�̝חr=�_yȽ�	��q��\�t���r��1+�8Ё��(��+������,a�{�X���\զ��ߎ5�8>�R�c��1���N�I��N�Ѫ<MN���D���8��.�����Шf��ǥęF�G/�!�<�̹�ǬK�6����y�
�Dպ�r�:ҍثs�֨|:��ZT�}2��-�B_ZF������Y��6!�ֹf��|g{m{fǼ����kRaN�"�n�T���f}��KZF��ֺ�����dW�����+M�)�{cm�T�7�wj�E��a?pVb߸K6
�%���u�;�u�~�Z�����-$ۉL�
7;��������u�#�g�Z9VLnt�a��+֣�T�G�s�b��c��hר��ԚZ�h�g�yç�}OU8�W�[8ȁݮZyY�e}������ރ5�V��j������U�q
�'$k�{|��N8���� N�d�����{N���z���V*�3&��j���h"QypȀ�)�]���1�l��?��{��ɤ�W�*�\U1������H�}^��XO�b�A;*��vY�V�?Z˭�fԤ���;����:I���Ѧ���V���CޫIF�ǙO�Lt]��\�
�_���a��5��Eu>��k�
ǚ��3Bj�>θ���>���J�~ϩ����k
��=L�șઝo�ǔ��|��򆖧*T|�K�Z���E}t�q�t[֮pZ_^4��'q���0��Y����G	)�
i��f��}��}��{�#��F��xb���1J�t�S+�� �{��'�h�]���������+B�t���H��`T�0����b3t\8��O����K҄�4���kw�zjD�qV�hlLsVk�Wt[~_1�B����'Zm�ȯ��;3M���y,u�yV_���8{�`���k1�Gg����ś�+�z9�ʍ�o�0�s6�N�7�ä%�z���5�BMw������r�Q��iP��\��S�q��2�� �C���Z���@��s5��aڡM����,���#�+�'�׊��:$',�?^�>ܪ���9w{���d��=���q�6����o���8�����i���U��{$�'���e��\/#{����1L��m��ð�q4S�~9ͩ[3�c092P!����ʵ7[xv-�y�Dc��k�Q�mV�3O�v��������-&��Yу ղK�����)��)��/?�z�*�щ	�_L���o������s�E\�I��ڒ8�r?�uB��XF�����J�Y�����6�te_�\�v�}5i�ت�3�YJs�p5��v51���Ho��=&	������N����,ګ�>��-v�w�T}�=)mڔ�>�$t@Ajw5-��y�|��HX�F�f����=��%n� ��z���4��[���s/-j���c�͌	��ֺm�M�F5�����g૓�/��w��n�E����WS���c����p\�S�ً�t<�/o:*��=&��v�>J���(}�b�pE���s��B�GH�Xo��l1�Kիxyy��n3�^��E�����c��_�s���N���ʹ_�.��W�Z����K�c�}]���\P�}/Z�k+�Ć
�_9�fvE]��wT�$�91ϰٍo��kj��s���<�vb��e*�&�=W�1ȟ���]-<�Ү͎�2 �Ē�5ym�Ѫo�1����_$]��c;#;?���c#6�rsp�k��i�4�-�ɵ�I��G�k�����1d�{V{5Y-k�
�`��<��)�mr�I�~Q�Be^�9�9:/�(> #*�p�p�<֋�\{eS���S�7lO'� z|�~����>3.�&"�q}6�x}���lpr��+�ڐ����Ne�U]:���gm����oNhVU�f���A���%��;>����䙵m���ck��]���S��?�Ty�漏ɷ���0��8@M�`�N��@ ��G�����{
H�9�h>KM6oV�賀����^c�����>�>a+�L|Bqр��$�������:�ɕ~uִ��9�Rآ����}�`��q���<��^K�ȴ�B��Tb7;�8�k�]'�%+��]��%�������wT�T\�'�e��L���E�J�4GD��phX����#�z �qn�{;�)qz�}�C
h=�Ɍm-)�v�Pr)��V�鑎Q���$��ȽRcG�x�枛��������k�4^�{�ve��|�_�'���"J���xj��F}^�CqV)}�M��rԛmL\ov�^�)N$���Vu����L��D��F��͜
�05]�r�����K(��|�υ���F��=�"�3��%��hi�8�ū��n���kKUp���P����ܣ�}G��.A���"�e�(,W�K� �����H�~�N�:�����S���Ee;��l��F�I�4�WO�y">��	��$| TF��yYe)�2�0т6$~3�]�I�յE��Z�o�~S��sũ��"���	���G�/W�p��}j�H��}m��~�Q�i�x/"��j�䨯e�Ϭ�.���)%F:����rk��֬�&��r���m�ĂP"h^�e�?�f}�|� L���M4Oymg
**�l�;�V�L����IeqZp�gX��%�l��)��47��}i�����4�,�S���>i�>m�>e��-���$���*D�hAk��g+��rh
�m��~d��M��rѕ�j�5�����L�55Uj�/n��P�%�\X׉�Ѳ6��'��/%NY�������E��=�~�`iڢww����L��W�|�B�j�_OR\1�P��G�����?�>�?����Q%3�S�2NB{���!��4q��Rо��[�3R:g�<�_�P%�~��������������b�~RK������A6��iD޺W�/�r�ѿ��%�F�W��3`��3�y�ݯՋ+1�
Sу�꓿n)��H��
չB����BS <��q�J������M����K��l4����I3h	��re״b�X�ۼ��ü�3�tU�ա=�,&/�з��.:��b���f���ѾA2aS)h�s ���C�J���Bű&��ا���"T�2A	
��i�-�4�-���zJ>_����m���9��'L���8��@�^��xk�i(% m���V�=b��jٲ�%�D-q��Ep���g������f5�Z��ĳL ^_�<|����,s.�R����Q�%;z����aht����ě�E[���5�K�K�W�s<���!r>�s���GV����o�]�v��fwC4{��\�w� cH��X ���Ĳ�Am8�{�<�(ThU���ڰ�����˭���7�;�r�x቎�%�Ez�����*vU���'Zv���aw�Gp���^ʆ�O��k����^�<��
T�D�_V�S�~}���{����)�j����K�:7M�1�5m �P�&��-�`�ok��rv~�"�!?��h�l�:���B8�­�/ʤҪ'��լ_�i	P��8���D�%Gb�L�&OZq-4?��3M��V��t�K����cW�E�
"ӗsiH޹ɶv�H�˱��c��^bɞ5iw$=o5R޼=��"{�bIa��*
�29���x#?2�(��;� "�t�M�nĈ(N����$������Uΰ���Qx� �f߿�oh7�V1ov����G�!��Ŗm)0�fS�E(�E�.Gp"�5��=;m4ڇ�c(Tq�s��t1�2���R������Ae|����ĭ�~��ms?p\���Ӱ�4V˛oq�r	����u�>Bˆ�~ey��k7}��7��0��@(��ߌLA�pf�?���2< o�P��gB��P�[�Io>������d��c0�̵�H{㸟��Q�W�n�_���e�n�5�5�9��Diw!��9R��SMM�ԣ��X>znfn���|�d�;Ϩt� �v3��n{ad�ɽ���.B���4�-,,�)}�}�V����R���G��&�Xz���-r}ru��"�2�����O�C*#�ڿ�S� � ����.�LS?�|�fzc��W��pe�]n��m�4OJ#��P&��ֺ��%?�����^����dKtNSIȂq��m4+#&oχu���C~��i�@��oF���|a�4���'ٷ�L��.�pf˘�mݯ��Y��u�7��b�s��.�'wYsp�(3&��)@1ނ���T2��P�C�̧�:˨����.ny?	������aϣ
c<��w��R�2����m��m��)O�����~X?G����]�#��+�|���%��������e�����}����o���[���ږ#X#tP��+ƫ�M�KmF]u�M������&z
8��&��6�]y黓�R{L��<.:�PM**]ˁP�ڽ؏�vC���r;�|C-�5o8�u��Z[|!��w��� ��ڧl�'�5���$�d��o�S�� 3ŝ�[��Ͳ�n�'�~Aj5NR�ʂ�x�<HA���W� ȧQ��]�w1^���IX�G�7��0Xզ��n��~󼖘:a_�
�Q�/W$���'�T�*�`T��x���u�g���͋p�:�߭.��Ŏj�����Sh��ҷ��e5�y�)��:�0n3)�O�
	_��J$�(�Z��_�����$LXd�$��5;�R0X c��m�&�23�7p�P� ʦ����e���"V���?��%�V б�L���5K��^�Z�ȕw���s�NRy�5A/�`�̭{�"fХ�H�v��ﯥ�J�j�9��r+9�7�ŒR~zN7=�C�,f 9򞻬%}��x+ܓ��D��65U���f�r���oxC�8�> �NE&�t�	#�<��|�g��X_/�ޣ5�M��	r�G�#vc.��ME�%ht��_�2-��N��|�Ԙ���\�,�:���Nl	-@�p�S��R��v	�
��� EF��� ���<�
����n�3E����WH��'ld���.#m���x�}�J<<��؂�O�/K�~jy����tP�_;0���L	���b@7����Ylӕ��<]���iSa�:V~���u��^�*��4א��B=�y�q���]9a@�F�в��{eܕ���%�7!2��J�:=�h�/_��D���u��x�h���G߈��Dו����N�Xo���(U�|f��VK &�7��%�IcN$͗K�p���x�"G�JO�v�s���Ş=K��Ƽ	\�sY�-���>����U\�;���,)JM�a��`��
xg����u�\~ $&��+.2��n�O4i��#4Ǭ!Y� |����7Z��d�3*6��!�o,�.���̕�� ����#Ϸ����̕bC����<0��6	��h�~�吻�/ۙ��I. �5��ȂzB�!�ky	��L���珺�@�V���I�#�B�3�_-����,>�?�������g6�zV�D��p��'�l�3hj��]k�T��i�W�4e�n�m~��|�Q��2���T�S�]~jX׫!T&���P��[�3��8]xk9'	�&(Z�m��0k�P�ԩ��o8��⫑��#��1�N��/�KT>��@7��#�)[)>�8#v�$�L���DPl�	�d?MEY����6�q���i|kԫJ�s	o��B��?'Fz�|u�x[[�Jh�9�
��oM���DT�� ��5��=��7���\��Xjm�.G���H�.�Z� ��#��)��	���z��1<N��hN���m*k��>yZ�P3:�wܦ�ޱ����͠º�}n��	]>pb%	�`�w��@ܝ��~��~�
֛Y�G���P���̳Q8�+��s�8�o�$v<=kW�9�Q~���b�n�x����Q^ z8Ʈ_/덈�.��u��N#�gxK����Ӌ��������ȷ�x� �d����ӿ�m��%�|��n'�qyK�h��A�n|Y?̜);��L�tX#��%8H)�W%L�fyS'P�s�odQ�|�eD+A*�ۀ=�[�������y��Z��}�������vD���� �� ���Xw�@Bޱ�p�����s�&'�._�B�&72LEZ�Vs���*�"�?B [ n�F��
4a �c��Л������?.��wj����Wc�;�Ŗ��r~\P̶�n~[>V���cR�I��R���� ;zPa����i,�.M�"���s��}4�x�)F��g��*Z�)u���);�E�r�kG�ͳ���Y&d���� �[(�������6�X@8M��ID��9'M"��+��G�s�H�9���s+��;눏o�[�� ���7G��*H��7l7d�S�y�����_�����*��vw;[=�(eNT����#y	+@����7O�� �� �����"T:�f`��Ҩ�2�ĨC*�N�0�/�kC��kna����D�Ȕ��d:",��z$6��'�t�q]�Kp�F:�j�(�:xd��v,tQ��f#�G�Z�k-$4��X�b���Z��daO����sT;FB	a1�^$ԣ'$����G�r�.b�v��mQe�ơ�e�<󏾻�S���Q��m�*/��J�4
�@%�3Y0|�O�T��5Tf�?�\�C����Z�"��ݩ�U�2;�	����s����ui�{:�Z���ɕ\��ʅ���u�-�
�����y�LMx+@�l8�=�E�Mx����Fj�j�����h����w����@��3���S�6T�@53���p��2�*y���K+�ۓ�*KH�$�@�0�)S�1����X��~*�	n�˪�{]��Q�9t.�g�V[�0��������j��۰7�O��\A�UPg�=_^�3��j�hDl$N��k���f��>�8
 Y�fZ���` `��I��t��0uўzr0i3�5��Y[*���>(�0�-���0�q"i��=|�Pц4#3��nW��c���gJ�L2;��\�I���P�>�y(Lƺ������V�qSۻ��0�a�`�r}�(#� Ʋs���g5p��k@l����g��X�n�"fٓ�'_���0���}M%�s[�y�����j��Թ���2R;�S4�{��HTlĨOΞx���Yx��6w�Z@t�Dv�aQT+)=���i֓�pC�%����8����D�����	b&\�=�l�U�ð@uܷ��uM@h�ܽ�Ǹ%M��g�����s^�@�mZ�_�yY.7�5lݼ�q����	��Y��M3;s�'�d�FN�/��s�ܢ7�T�A9O}�&
���\�@]�d7��bsR��w�9�C��&i�݇O��.4���VH��L2T�~ �fY��\�2���L�&�R=fL$��_��|��w�-�ԡ�(�������v��Q7��`�5́L3߅�@�f`�1&^�#S�x�w���a4��m�	�{�����<K��Xw��מsR%&��7�w%��u:�tXF?wn�Sҍ�J�aC70�A��͆f�hDE�<�����G���|�/~SI�E�l�U�K�u�*q��m�>*� ����CQbu��u�I3�C#�N`F��Љ����Dm�sм��( ����~ �o(����W*���\X�t2���4�tQ���kb��6gl�Z ������[h�*���_�H�Du�e�&�% 	�:��w���M��~��OԏtƔ˙���_��x���]� ��=�@̱�hȄP�t���5�I��{],@�����U�q�k�`k���G��Tx>u���R�+��R�.��l�����EB�?17j����om^kdRI�T�k0fQ0��5>���@yl��e�1�V���1")����v��K�h'���TW�|ŐG�w�XΩ�`ϑ�2�j�?�JMx5�
=Ӷvʭ\:�N:������g�|�7�H ޴n�u8�p���7x]� �^# �l`�^���;(���o��'�Or���%���pVj�-~�m�7h�{��M|�1|Rh�R[��`xi�L�Ӡ�4hC�=2�F������֐�֜�~avi�d`G� ��H!x�$g>���>�唋�
s�/���
��djMQMؓ���&��9�lfi	9�����DKrݜk��]ǥ*�0��ubhw�E	�i���*�p�&K`X�3PI,"=��?C��dŌˤnn�ܣ(t
n�� ���aKm5 4�q]jW��K�aM�|�1�7  ZPF ��|~��5g̻WB��P�����}�≘���O|F\_Z'�Y��:�(�a,"ah�5	;�������_��� C*ҭ�`#��$���?�c�[��R!~�hS>�=���M�f�����(�	[�z�/��dL:���� U�g�|e�`�ª��(W=�Ђ�r�둎4 �����/VuA���Z0��U��P��J��Ե�@P��砡>e��W�T���tZݫ����z��Q��I'�=�I.�ɋ�Ϝ�RNh�]��;�����P��g��l��������3��7¸M��l�#��eE��^H����!M���'s>��6,v��uߢDE����O a.
-��'sR�M�Ō�x�i[P��|�G�e�b�tC��4B�&~䪗r/�pR[�q���]�[?�bƕ<�$��+���5��:�Dy
��w-�֛K\t�������s��:�ˡ��w%j��?�!�s��G���ں/I�Z�`%��0�f5^L�LhG�f�f5�� �o�y����j�A��4h���x	Y� =F�2���q$��hK�>T;I (dsN�3C{M���%� $O7m�{��2������p�S�4C���J�	��Az�!�+��Ǯ>ZA��kBk�p`�@���La��T`�r�L�qC��@�rĔ=���QVd��׊����G+ �<Ǿ�۝��;������JLK�`X�j�= �h�(�d�{�@��s��#/O! 9ۡ����C�r�l�_<�����g�0z�&]�l�Ǆ� �%�7Y|+.�T!�TU����~����NL\6_<Zu|�R���r�r�_�퀷_֓�'�z�2׶�V�1��L�U.7\��������b[�tȅi����sL�;G�u,|ɢv�2{U�vOL�e�<���$_�}��U�%�C/@��� 5�2��ÇOⳅ�#b��^S%�
?L�o�h|��A�Y<4�,,XUU���m	���04�5��c�Ix��|�\׸*/Mw	�5ι~c�|o�� )��·��)F�&����o�+:fїO����w̢{$��ZR
B��[���+ܯ|�t��ظ�m⽃#��J�	�͒����و��j]b�	�"�5�N�G	nu�������v�<����D���]�����*6�]�70�|��W_a�w8_�����(���V]��ݩS����nvdI$�|���m/M�E�o��y���t���}����J��0��[6)�{`ĸ��0-��F7?>����c�ASQY����3z'�{�3V���#��^�8lk5�7gh���{AE�����V��8b�K'ݓ�����{]w����T>�#��L:�
¿�U����4gO�$V�8�\"dciJ#N華;��ӕ߹�T��;$�Tn�i��ԗ�l���9Κ�gۜ����|Y�1�C��h�^�S�4�dU�C����ۊ���%���m����@��7 ������X5�)^��#t�1�B{ř�D���g�V��3��l=Zc��'����ԕJm��N��m�U��u�=�tAo��g��_Eq�H�gX�����j��tu����8�ؓi�=2��%�;���t�z>e:5�n�L�Y����j��*�5�RL�3�ڟ����g���|={������%_�r��j�	�M�x&s��}pM�ʧ�֕Q�=��˳�\�x十͏�rW�',,����U
�̳AG�OU7ߟ�u�]��b��<2��E,��l'�lf���췌�n��F���ò�y%L�&�H�e�3�OT�i*)�������'�f��o�G��߅V��H	�O��t�sa�FfN�fZ6�ę���J�=G�q[ �s����)|)��]��K ��S�<�W�؝u@��N݅����m�%��ʱ�4c�^�[Zh[g; <_]6-�}�9ݤ��N���-����h�(w�7�y�zxU�~�'���o�yԴ�m��A���|^�<��Fџ��E�[�'T�W��U�-��W+,+��ˈ)�k�{�e�7�:î������6�Q[�$��{��@�J̆G{b��-ĵ���Ŀ�ߌx�t
�3�y�s3�g5�Ry��J��Pw�{=�p�th�WO*��H_�{����'����e�$��͏������M���h&zS��Kz����2���uU~{���`�N�ML.m�:|U�g?�A��������
l�/T�1�h*鵷�Րcfӑ����g'҂��N����5�����2w3��"�ThF�]�������T�;S��u�a�&����f=��V�,��)���rV���P}K{��~�`��E��#��9�O��:Έ;�Qe���l}wr|D募��=M��_W ���$�9���ad9��cs�#��8�����S0⯆\�\��ȋ�9]Ǟ�bj'�X�����w*�`w��Cd�Wu��PZ��畭����]�<j�n���)(0����_�'�̰T`{x���5S��v�L%�T�ۦ�</���̥mx���e�a���N�)���-lrm�$�^�H��T�-^�z%D���ǿ��w/��>V�{�t����L�w��BT�C�������/��SQ=!0P��d0_�~y��0u��p�M{E���5:Q��%:QCt���V��^�GQ�wV�{���,+���x���~�����{�k����ϵ�0��m5� ��D&Ja��=��Y�TT�Sx�Y��z�
~ω�9��t�!w��C�������,��������JJ�/��V*#�����-d����ǵ�ֶ*W��7�ҁ#�{��u��%2e^�q
�gW��'�5��Ƭ7�J����+������4��?�g��^Y� z����@M���3����6�`�)z5��9&����
��m�6��G�*�NO�󂤣E�M�K���;p:��Ԋ���[�e��q4�x����>ə\�Y��@��v��,�\H�<�e�!>���=���C=R�V�+��"�mzC���.�ّ�;ZS�V�o}�$m��pV��A8D� �9N'F�Oz�e
$��Hw�~�I1��'��v�H�J]V�|�C]����::J��q�V�����	4|��L�)��J��:M�0� ޟ%�=�nɚNJ��|�ְE��J�?>�*�LS1�M�.�y���(��E����C%�4;7�;B߭�&���:ۋ)�0Y�K��a��ގm�k���~�ݫ���?������a�����#qA�K¹,�[�\��� :�9���#��� ����M��̀�[͎��t�{��o�Î�R>Г����ҹ �R-���tK���R0�ߺ���w�YA9:Vs����5�Q�7mM�^&||zcTk6:�a��q�LO�4*�b��W�v�R�<]W=+̹K��M7('�!��Li��z��Y�2�`�T�t�/�t�̑�z��iV)��"����2;Y i�ÿG`�FI'PX��J�����=r�u4������&Ǯ�cBLL�
X�g�Y>L/=k��`:���'�'HN�����y%�ǫ�@�m_�8'm����e84m�Ͷ�/���V`m��I�<�]�l`W�+�e}��2p��Q9�N�=�����<0�w�Kϊ�����3\$	�R���/��)�BG��<^=`}�6? �Dz����+�ط���o����/P������3t;�XТ҇�W�[�k?��-�I'X����9��8s_�|��g��sݤ���t�a�]a���{����<�xF_p!�D���b� �5��?�ը3�����6>�H���?9��_�Vכ�ݧ�2/���qR~�?-5Ld�hh�=��k:�Q���#)m	��8�C�	��G![���h��(_\�Mk��ݧ��K��3X�?K:��~��,3+\�5�V�q�0P�J߈����d�ȴ�tO}�۩*����ܱ1����Y묐�D�j뷯]�!��8�*d<r8�>d��G��/���I�Lm �R/���w�Cע��7�.9�b��#�������:�X� ����������+_� )��9��A�)��l9�_�a;����*@iS���2����T`T����X���kR�q��Cic�e;��|� ��1_������)_��!4��è����)濽��9����:=7��s�1��a�y�	��9���n+�G�M���E�5��;��(����m�|��8�`i�5�Nk�*��4�
 _�M�	�>���[�a��t̍������ۉ��b|�0e��G"�\Z���a�R-���z�<+H0^@v�e0~�r|dT��q��˹�����aR�kࠤF������>�DpΔ� W��f'��"1�9$�q�ҲG�����3�����3d�SR���UQ���2��A�1dboS�X5���FbS���](�ȁ"�� +��.���ϳ�|���r��k�f��>�CF�+�ЭP"+����tq�Y�-_�*рY�5�?l,���)�h�c�U��ẏ�3��u�&��o=���B产��9�#'&�:l�M���u83�RQ�]V!���h=�4�վb��Y��V_�����^�=4Y/���j7�dK/�f8y�tB��D�#=�� � I��DC����u��O����������t4�j�(i�o��s�=��k��xJ�cj$�W�h�N/�xP6s@��z�q����^Ced�Zg�F�(U%�}``��2���a�[U��#F7�Z���=��ŚNb鞹;cQo��*8"�ޢ��V�(��t�ݙ�PN�VJ��d�y��%����Y�2����M���[��U���_=�����ѺCF�����u#H4C��������Rn���H��e�yGf���H`ml4�ƀ~a L�w��_�\w���D�K�/֤�֋�O��N��l����2��k�s�y?I.s�ek��?�ʾ�I"n��5��q"dn�u$h�z�i��o����w�rms���s]ANSD� ���a�������q��/[m�P����}����ZW?`z���WU���%X��~Ne�y�!I8�y�.�JƜbM��+��妌P��l�s��'*�[ُ��f��2��rM�uuS��׾	 r��s��
�)��PpA�|b���,�Q#]����M��\qC��g|?@?�����;g�l�W6�B�،�W����"}O�[��U���b�(CĜ�;_=�v��T���8�M�	B��2�ݰ�Y�_����K����8
-���m�_����.�奐��s8�G��E�1��z�υ�8#q�S١{c���ϗʝp�ҍ���p2o�I�f~�[�(�����`�%�e
)V3�<>(ǉa�l�	���SH�Xͱ�^��G������7�W�W"S����[!��#ް;p�H����L9�=�;����)!6M���3��suRL��^�r�&�F|!�@J|pEsx�؟�IB�h [�I^CBv��E{뷻z[��塅 �@Et�����w<:%6����'����"܌萸a�d%m��������Pc��B���P�n֨
���ʗ�f���Ǐ0tvf����N�Fϥ�俆�Z���Շn�p9�&���C�_��|�H?�A�]�Ob{٫5&,�����*.4P��s�0�*W!
qwG=�#Ry/������7�%K�����!��?�~U~�xp�#����*��齊uE\*&����Ё��C�ҭw�԰3J��g�����i(����bn�Zy#D?HӅ�|����D���om�.D��X&˚�mH��U�>X�=�+.Gw:��<K�8���)�w�U��W��5�J*���+'��8w	����S���6&��P�v������J�����S�Ĥy�eb��א"/�TV�.׾�9���Y~���E�}���ܖI�:۲4��<� n�8��MHպ�0]s���Q�Ϧ����v�|���E~������P(T~x���t�;�TBE�n�@�6o��Tv#6�ԥ�z�����QJ AH��.�C"�2�-��S\������\HR.��)�#���o�6�#{�`�e���c��=�����X3�@px�Pt@D�Ǎ�.�.b���soұ�*��@ݛ	�K�Ƹu�mA��������X��qt?Ӆ�Oށ@���/W�>�A�?�^�t� D�D���)=�Ó��T}kL$��ާQ&#�ZVs��Ѷ's��܉��Sw�MS֥g\-�?A�._��!ߑ���gP1��S��|�+�Ӗt l���M�$��/AA�ö�L�6�	1���Wm���U#x�ˀl�
�2;��@�C�S��)�.7����R��w��W��������@m?���&�o� z�F��B/j��k}:by�T, O�y�]W<�1��k��$j�s"F�'���sl=t�#a�޸����
����4�M�E�	�n=�`sQ\Z���tH�3n|g���[> DCP�l�
_QM����_�dB^��6��ɉ�z��aelv�"m�SCH��+M�N�K�np��T4��"�����O_����ASL����<H���#!�A��jTn��dP�!���4N����^��{M_�Lͫ�{����N7o�a�)��*z蛎	���`,>5x~��!�@�6���:�Z޾<v�I�[�
h7���,\*��N�yUۚkF�o��� �9�ٹL�u�o\���x���7�c�����P!�,�U���W�g�C}9�N�g��+׬L��FT/$𓈕L�@{��v7ӓ���v�[d�0�ǎ.�����:,bl��z
�X�0i9N�,�U�����@a��DX�@d��� p'c%~X�n[|�h#���Cl�{������A������jvZ��*��EW���԰</�[�3�=d������,Om�zA��j���E~Q?D�s|���dl:Ǧ�p�Na�k��P�������x!~@!\�����Q�}�����W�~?�!�����1 	z�R"=�3�$nZP�A�d�*�ѯ@��ۆT󭛖��h_�c,��o�(��|��r��r^Ώ7��0^�}���bO�1�B�b�	k4!0L�D#&����n���=��D�j�!='l�%�y�(F��2�=��U����5��{���N΋-ז:ˑ+�'��j�{#��(��0���	����E�g&���i���?p�gaT�DZ(�y������5��%��Q	v��z������x�������-P8�-r�pgU<o�h}�є-�r�,�VF�`n�R�^J:/�Ĵ��*q؈��m�٧�jj�bKΒ���O��I~!Eek�<J+R��*��|Z��/7��,�����"�('�tT�ʌ�����gA����OWq��=-}��\]�!�&�([���^G��
GM�/��־��3z��Zt��ȱ8q;�i�5T�����u=��A��O�O��]����ⱁ�e��������9�rL�����H��Ʀ��+1~I �n��CS�'Fg/Y~�s=�ػفZ�"����΅ḃP����X����&�8�_�K�ח[?&utej�Yގq ���W>-3K#P��dϦR��]���]�ժ5�J��a�a�����!#���!��q�S�F	fye���u��@F���-(J�0��+ܱ�\ԛO���XL��&������.@G,Y�u�[���94�<�C!\��h)�]p�s�	��u�4_��o�2�[��_�+�)1.�o�,S��5Z���D$c�=��}{�oȟ<���o1	���&�͍ն4�4���W$��x{a�v�[�OXڻa�"K�����[BCM�4(۠?�!����}M���/�/-�)�C?��� ���6���j`sh�G�-җJ�_�fo����z,'<�
��\�$�Hг�	'����mcx�bmtY�y��`�_���-qk�p���z/��O�"�!~�G8����.S���e�U�����Ĵ��L��ӿVC4�:uU%�+���#�^vf���]x�8#�ɥ4��m��?~⯘�ts���䯍aH|+���bV�98��
���?E5�����d4����_��ɜ�b�?�j
�e�B�;��,����:^�mL뚷��p�j-�C��6��B��`N�d��|������(.�H"PFmR|�ֶz�a{(D)_yG����{"C��k�mڛ<��l5�&�NKBΫ4���,c���WN4�����G#�\n�0�տ:�=�*mΥ�����?_���2�����ML��,�Q#1�jU��֐،�~�~z_�Սy����6�o�)�E��.�v<�h�zZ�����޸�YSn�>J+�}9���O��}}��w���ɀ?7�oS-rM}�#H��%JP6X;��&�:	=�δ*.I��`�i�d�2N�.bH;���c:[�1��k�v��`��⑲u9q��#h��V$%�o�i	�4�e#��m�;|\*`ٳ�e�e�a?Hc|Tý���%p=�/ ��Zp��'ް���΋�#c�=��8O)���{�	݅�ԗ�o�a�Jes%/fef����'�]�m���Ǯ���mY��s��6'!�a�$�I�oHd
�V2�O[K6��|���h����Sh�iş=Y'Ɩ�f�<�22�|�G-�����?Ά�f��%����!�*A��U�{V��ey~�vq�����GDG(�~Wo�9��F�����j� Y�?�v8�cK�L��7�L�6qoY�.�j��I���^�t
י�s���X�À��2�V=��B(`��v&|��r�1ϫ�n+�{]���
�r�b�u<U�>I̘��Ѧ�������l)�tD����ٗ��s��:`ߝ�JMaIPkcn������Oρ�E�R�dt0�c�S9��غ��9eA�P��c�҇�u��YB;NB��`�YOM�]�K�i����'�ϼ�^��I�b=B�������8�im��[��	�颂r����r{Ͻ��J�@��8ĸ������v�5�e58�۶Pa��t�G-R�x.R���*N��Ө�ǿM5�q�jѹ��,J���;WeGC,�gt��H�ǉ���Q�\�/�2p/�����[&�:?��(��ړ������n�%
���B��I+����K;�靺-��\Ƣ���y�v�s���Mr��������X7e����9*������rc��W����(����~�^�2��qqJ
4��o쓇v7�õ��E��j��D�2r����U���Ï_��I�?�B�jE e[��Y�+��#>6OZU�B	��
��a���d^�`�/�ۺ@���{}aL_����O�����_l��G�+���YO����λ�'u�dC�����)9i��i�u�7N��U�G���%p�?�~ׅ��Z����]I�(�y�PPC���)�%�mlm���u�ͣG���.�e1-����zd�\X�^��c����:��a뿞���@�+�p�x�����*w��Ԍ+l�e2�F4P2���@LJBAn0����T׎������N�=��h�R�h�_����s���QE;��S!��3�/��Ϫ��փJ{�s�|��Y=�:����^V˱ʦ-2��~�Ky��Q��Dlg���Uv%8`[��o�e=y�Wa~w�g4hɸ� �3��5�/�qT6a!��a��p����"z���W�OL��*"Y���w.J���^�Hv��%a��$d��ě��e �_'�!ߜzN"-}��T�{Y�D*Tx'H��\�3/&�)_���[��L�^\OtD:���.?����^�q�p�17���U�X�8arüOT�l���& �4��miR�����[�9C/��>�8��r0��ꇡӯTN���o5��C��ױ���T1.��*{l����6�ۤ�п�s�en�wK�m`t����d�o��Y�����ܟf���Os�j\ݫz@���~�7�w�BIE�Y�y?Ƕ��=�ION&�0EG���}�GG�M��e���;*A''`��ޭw���`����'л�D��2�0-�,���_ndO���f���;���4����嘆��gq ������P��9&�P��I7�̫ˤ�*�>\�|0cgV]����8`����^�4g�ٲ>���~������ER36�6�&G�d ofe�6���L�oR=m��L/��!B�N�K�۷��T�y��o�`�Bf��Ns���l���r;��,�$%w8��`��ڌR�����hl��������(O+�c�i#�F����������/<����V�{�_9r�K�70a�~�p���˧1mb��|�se�0jU?{�xo�Yc�7'�X�4	W�B�n��\\cDp�c^9IL��q���E��p`�!�����,�4W���*�`�w�Y��6["4��,ö�J]e�A�؟|� e�$�m�1�gۋ�r J;�s���9_�ߢ��_"W�@��wUp3o���Uk@Ė#�g+Rb�>+��-_����:a��_�Դ�!�* jmȚ��5I|!�ICT;0|���Dy�
�oV#���@7��q�b�5|4,t"9���Wv8��ĥgz�bY{�뽁����M bJ\�CV�����А�訤O������Ы�X�T�w���ȓNX����S��4���Br1ǒg6K.�N�O�����W��1�n��L���&BQ���RO�%=?��5
2[��g�ldh��b&}���f?v��{1��v�Zw��u�hs��bF27VO;ω4��X�G�]�KT���D�}.���/��0I����`'i:j��sC{�W�����c�%����+k+U�Ob&g4�Se���/��A�8�������QA�K��2�.	'�pjBrb拟�p�L�N��gp<��B���Zeyۄ�v��t���RO�Q}
F��+'Y�g�'��F���N��X��W�D68
�;J��9V�"?�?�"��Yw��p ��txh�4u��E���Ds�����K����V���(� ��XϏ��ݪ��Y\��f�bï���'
��ܷ���B⪣�$Y]�]���0jf�z�d.�%:c��Q���.�>T�-L����,}��� N���.�bn�7���]'���v��7���ީ'���Â �*����bR���}����#����R�UG�,��b�1��#��N� `-��}i�t�u<�ܲ�.��0$Q�����y6���C׿����g�ge�XC�	�4�c�E�����&_-��-�D���5W�F�1��w�;"�ۢ�𡎤Q\7����йd��_HSk�|�_��U7g�!�[d*.7m��&��;p�.P
��r?6a�/�A;��R��l�S�A��-�tD�p�U*f��C��wY`�>�fN�H̰Rll�~�o�'��3ko��O͛c�w;��"�������x�Ɔ�D ���1u�����տ�(C����'ۅZ58���Ż��k�u���-𡒻��bt@�����'2��B��FF��������R����x,f��_;��z'O���W�!�汎��K�:����7��(�}�&�ŭ����wsx`����iDP�[ 슺��/c��Z�e����y��a�D�>���z�o5se<�o֊�'����-�������Y�)�p������߮�8�Gg�pe$ݛ��^[�[�Mw���|���>_�޹��'��[�]M��/~��G���d�"M�4��5Or��OV(���=[�D�0_Y���m�~�`����*�T��1�lX�.0�prX(<�^�������Htu�=	�v�uRY��E�0
'�G�5��?O0}��[��jJ�5"&�P~�F:J�G.a�?l,�����jk�A�� Ir;�s&y�й�ɾ���_ù[��t9�:�w"=�}/��RăT®�"��_���g5»���-xᯁ�1�h��O]��EBy�<�X�
L;�{:�4Z�H�n{���E�F�GBM4LvA����y0ܩ���d�C�T�贐/�bYē���L�	nu�5�Mپ��%@�M%F.����׾tl��r��S�j�0��+��~8�$em�y!w͕��`*���%�&=�����A�B����؛��jU(����ׇ��T���]ӿ8�3��;�pz�ss��OP6�O[�2����tLz�J;�?7 ����io����[{�O@������m��wS��~}ie!�/O|�1���gu�� �,X��\\�IŒg�O9F4;�ǿ�d�@J���SPބ��W�zx1L�m�7��Ɛ4�;>�b�J�=s�̿���ҝ&��eP�q�o|R�K�*)a���nC�����wY�����T;N4gj�a%>�sLh�t�=5���)M5��|��B8��f���h,2e��k�O��+�l
��Y����Ox��fmŦ���x�W��'bS+��J)s�#~�`��}ԃN2"�Ǜ�ő�E�d&�kH�x)U�nL���Y����Or3���C�/�,��Z���T!`�~�P��R+P�oM�����¢Uw��E�3R��U�)~�<1���Ga/���9\��weQ&�~�����E�k;�X��Xn\�).��J>^��X	?�LXM�� t��iӘO�œ�����{Y (���n��CӘ���w	��RE��c���c���s�o\�D�4�m���w�!���&���Ӛ'�M�L��UU俻�@�����_�a�F�#��ӫמ�Ŷ�πՋ,�!��4t,e�q_@s�M�4 ��+)}/�	�u�9�!��̾���A(:JR_�;�۫���=0 ��"}SJ���Qc�6�BJIs��+��� �S�«�^{��B�=z=�uq��l��<ŠA}_0�%���Ì�;�)��z.I8yǌTlZL�,'��ȁ,�3G��ע¸vj��<�I�����v�y����sB%բ:1e�@�@Q���g�'�U6Dh	E�Ov�A��1�O-Ͻ�兺$��c#�.��c!M��'��K���ʸc�+&����zK�j�I	X�6@gR=<���_��h}����^��X��hw�"pN�i��:}����qhڀ++�;BP4���i^��*�}n=�O��1鲡K�Ew��GG�h��6@�f�i�:�]�s�^�\�RJ�4�²s�5�E�A�f].EWen�3�#������8]R�R�9��KT�:��PZ�`1�h����wO���B��-U�(��l�Y��6�֥u�S�	?��y��_��n��{e=j�4�fc,�Y<;-�8�,�[�'����d#2ׂ���=�/�e�v<�o��X��8���)��W6j�O��s:�P�lg2���%���b���מk��x�|��Q�A��Mz��m~R}-���)ب��{��揝/`�%�׈8�ܣ_�8����<L|��W?Kp����*#b���Mc�y䒆 -p�� 5��`��uoK��T��034dHZAs�p �
J)���'�����O.Ȟ��MV�%��9F#_��J�r��{Q��Q���w�^XZmh��֚�ߑ�\��������6.���	�c�1G/�����=[�e�p���Ad�Q���{E��R���h�й��3�&��j��d1�`U��'-���G��z� -��C�/[����5�m�{�r{���ϕ�Ir�\C`z,�x��,�$W|�;)z~C	W��v�{_�ycx�>�D�_)����=86����,�;�xFAp6{W��F���]q��ࢱGYid��A�,E"ˇ^,�-�)�w �7ɏ�k���$�B�'���Bs�#3��Y�_҉���:�f-yv�`�����$�Na�*�:g��r��pN��������Y֤����b�L�h�P}-�����y�c�aRe�?��Wo�[]����ZS�����0g=ʁ6G�PK�K F�=%v3�,��HKCŊ�O�y�|2Ԡ7� ��8��>K*^L�+Q�����ʵ��'}�J�|cQ18��<n��bښ�
�{8L��|���|[��މ��p�֙V#y�5���&ACҮ�!��_�ŋ�	W��yVd�4{�u�aD�Lh�T��:��96Q��Ю��'� Նl(�V7�%�n��-�Vz�#�zX5@A�������ӦV���p	�!J��d����	%2^v�}mlQ���Nl8(�(��� @�Nd���;W1��k���O͟/����u��t�B��s�g��1u$a-�����o��v�0�8ZZn�I�ȪL ��}��+Z��d�ϗ�5��H<�yc��yiY�����5{&�{ޭ^�nD�]6[���W�q"Q9v���ٿ&���G�_P���"�ڎ��E���h���}mk�b���TYQ�#V�[�ƀ��W�O���_x���v�BK"�-#�>@�x�W���;�%;�@B�1B?a��)���_�������s �9��ƌ���9�Y^�������K��z�4����h:���B�?�%͕�ȁ�,{63��H�D2VK�	���1�td>�ybAz��'����x99��N"vjP=T��?�H��[Z�Hg!g��L�Q61=�������b^��.�	<nk���XRZW2n�$E����LW�ӫl~H�crJ���WQ��x[���Tel�j��	���9S*�����*Zz	R��8�/�pl�����%%�W�֜���\�F锂Q�q���2�d�k�4v+)h�����y� m���Nk�����&) NE�ӎ�����S�X�x��BȻ?�]Ε?7;q�3�<�gIm-� F&-�(��ݫǽ��$�@�?X��,���s�$�kt��j������d��_FD�R>_*絊����Z�޾-���2U�h�dN�Ҁ?z%��K����ٵͪ��Rj v�l�9�ߵ5;���p�1�����o�`K>5����g-�H�ITrLQa�9�I������o_�wϗ�<�mX�	zx<uIO�XÝ�����I&����1Ԙ�k�G�%
x�t�V�R�z�x�����N�~2�� �g�߮ʻY�Z��CǾ��j}�����6j/�ʊƭv&`�it��q蝜BT�s�<?�w�x�b�{��7�> ���}�Mw�6����0r�W��h���g�[5>%�*Z�EKd�kF��7P~��5.J|:�F�x��$����>�|�]Aw�w:�d���Ŀ�����F��<S��sL��W��n<�f�(��/ߋ�g�pP)v���i^�Y.K ���i��g�!u�UD;��/�ұ� �g�
$=�㇈[a��B��VX���S�x�y����m{�H+t<d��~� `�G)j����d�U�@������wp�F5n��pW����s���o������h|j�:�of��$��t|�<~���Az�5�k�vcWU�q_Ѡ��l^8��kg#�n3�5�к���2s�_�����r;7�!֨�uPO���'RQ=�����������i�m��$���ڍ����v���=�����u����M���#���v�agd����45P]FCp��3?�\�&?�p�-�+o����r��s��7�{��pPn���Zc���g�V.��/ǜ�#3��(�N���}h\��[����3>��x'���f����LHX��k�:2<p���%c�c�TO8����|	�ahA1�V�� ؼK]���v1�ی�X���~}���k�x|+�E)(��G}N�H��75�T�n:d�눕�h �n�D�G�V�gmc��!4�v3�>�l���"�>nB��v:I��$����>����Bi\���.������]1k�F�V���ѺT�zB��tY�P�>b�������:9����}*b ��;iY�9�1wwm��QrƮi�c�5?�Vl/��I�0��E�[#���-=^������_y��x���
 +M�J�-	�
���'X�e���3�?/�z��`�
G޿Tg4��=��үO	��db
�Ek�K�C���8�������黭����n*����Ĺ?ƿ�6TF.?�P�4}{�K��yhJ�{,o�E%���r;�wO�Y�hl�v�$r^	ډ��Ɉ�y �.�
�#��2��̚�\��҈��'��7��vV���0��ڤ�����* K¹b�+�w��7�][q\'g�)�A��ޫ�)��T$�=b� �۔.��q4QU�3�0X�p�E�P<s����&圹`����� Du�Lv�M5�)�V���=n�q:>i�gW��ՅU(���Bf���~̭i��%)Q��;�@)�B���|��k���O�Fɻ`�I��V�S�Fo�������y�G��!��L�C�5���o����G~�r?,8��K!tTG�G�8���Z��(��̖=�|x�lG��y�#�R]Bv�G��WFb/a!�yQ?�V*�����n��95�A �GS��j��w�3��r�viü���߈^��g��#$τ�Z�י$�٭� G[-��:a�r��3�����&�W�@���Γ?����qS���k�>�������֣th�����D=�%�ɢ@p���֥L�У��R_��q����E&�o@n��BOԏ����'�?"I�`&쇪�_������\�v1�H[Ӵ�8	ƜGPWh�K��`+P�\
g���Vx���~"�lܦ-P��ݺv���LB��@��~�$*���)F��	=��#�rb-�1Ѧ�
?Ͳ�^k�����u�7��XG="	�;z�DЛ�
pq�h�f����V����_�}��ߊ;Gǭ/8J%�!8�-^��A*��~�Z٧+��|Գ��gԒQ�ł6I2�Ж�$ž��4Nd�����I��������sܔP�k����<_1�`(�U�7���@8�Xߛ���V��8���e������o���Ï�oi���_D�i?1*t�KYk�W�v?���� ��>���,�ԣ�B�uݪ��s�2�o����S�,������6ŷ�e����*�97�D���g���֪��i��xT�T���c;�!ז�_	�MB�@�	�_Й�$����Q}��JH�ۖІ2ⓥ��K�c�;m�)csO�Y�u���;�2��>��2��N?�B��ZeQ�<ǭ�r K��U|����6��v����Ye��ſ�p ��9C;�R�k�����n��EI�]h�b�pb����?�16�����l�����P�ۛ^p ~"�HU��z�r��K�w����l<�ol��6Uy�X�SSj��)5t1/��I��.�N�S�.���3���/㼩�?�~���L�l<!_k�x�F���k�ppI�9iQ,�)N�v��˾�٪$7��9�);������NHJbs��cp;?��g~,)����F�j�mG�<\�2fv����+�*�v��c� ������'�n�j���l|�d�T�G3�ҧ#}VI�$��&�K�l׋F i(n��\lh�  0�\L�JQ\KD���w�U�>�yNNN�O��k��`�~�����Х��Vƕ2��6t�Q�N�~�l���gCw|$	�NO�:�'i	8�u��A^��Gѽ���DL�.�w$ *�4sw1>/�r�-�L��G��>:���:o��~���@-h�뚸^[92�a蟭E���m�C����U�`�fHj�7t�Pd�)��@�<Yw�Q7��	 �'B�>�Qv�9�ʷQ�7�<д{�U�z��/(2��ʼ��?0$?E�7�Vcm��|V���ۃ�"j���0��	a�\ E�|��1IK�r���d����h���j�m� �f ;OY��Sf@Q��vj�H߷��a ��(f�Z�g]��}+&���N��%!Z��t��`-���2N��t��#�f��_=�fq�̣��zrώs����|M�n �L46ن�L�t����T���Ye�&����ʀ`i����{�!e<D�&�^6�.�]�"���� z`蹅eÂ�r�z��ѵ�E���A߆k�j����kp���X����c������d���2��{��0���@'�q�M���/g�L�2>P�g���<zK�%��춋��($
��Cf^�X��<ۣ���u��G��cZ�MZ�[Ϗ�z��h ~^�z;1�Y���F���{U���x��*̯_T����|j�_0�D5��;b�>'�h�,s��������p���w�����+�i�[7!����|廛!�]�j�ޒ�s�����ͷ���̟4P�^}(�ܴT�7ݬ��!A�I��,����N) �k���%f�A�G9^�zT�ҁy~������u����:���>�k�1�0֠���1���yv�JTC���IeDS��xVo�f-Z����BX�����2�����'iF���s��|ѧ5?r.�2~�/Ap�1�~��=H'�u`�ze&���U�r��C},�����IV6�y�M��f)���w�fDY���2���EF�����wE�v�Q��Ժ��k�����9����*G؉�b$G+U�yρY �(;�D��D8� ��G��O֎�����X>����k��7Z�kFj�hcӅ����S�>,R�d������2��m߷�ye�ks�zk�;��c���E��T,Fx�.�?.��9�:�=������ad����u���9C@[�B�g�ސ���*�������J���@��9���5X+���.D�v���)��g^����e��������W©�'����O[38�5�hK��ZCr�1�����3�40�B$�6�a������#�% �\��\��eM�yk��a�ge�w
8u\A1ډ>�sV.��V�g�)���=.�9��.�/'�B��)� )(�J��\�/9ߵ���*�7�B��!��w���ĝ���J~���0 �l�5�Rc��F�@�M���V9/�a�ٲ��U�)�����=�~^��Ë��X��aC|�����N'g�� ��ؗHmuWݞuYd���ϞFy���^�$���{�vݯϖ��#���zP������������@���F&���))Ο�u��+��]��!G�cwE��
/9k*$�[k+�E�j�u57��_�s�Q� �(��ׄʓ������p��������o�/coF��JJ
�E�
�S�>��оߝnr/�>!!�L�1����t�>�\A��@֚� i�L�3�b������Vq15�P�}��,oF}|�fǔ4Qw��#��k����bnZ[���L}4Ҍ*�a�B~���V���Do�\��OqeƔ��Ӽ����|��ײZ|}��J�Ƨ�(����7���s���7�ᘭU6��i�!�v48���׻�O���uh�´�A��3�64�F��A��C�	���N��o|�����^�k����9�Z��x1�OQ�[�.�Xk(A����,e��]֌F'�[�ÝbS/�#�?��*��}D�"eЈ��H�tyQ@�;�E:�NE��.�J��E������ ����׺��������}���=�#DX~L6�Ng�eY�K���B�j ϯ�6����I/�\2~�|�cp�j�/�ܝ����-z�vIm&#�{7��sWR��82��IFq�,���\�ZJ��Ӷn� u�q�w!����!�)îO�M���JJ�8Bx��H�aC\�Q5��%U�$�Ga���<�[XIg��J!t���y�<�pzvT[,�^���4�T���z��j�$���d����!H���R�9��N,t5�o�c���3�����KɳMd16��P�p����>7�����lӛ�N�<�28���H���N'��_�Q-�?2��u�f�y�x�9�\�iB��У-//հ���|����/Oy�t�4ڗ��Bfre������0�l��}$�\2-gh|�%��荆	�0-���j'}~{�b|{.?�a�	_q�ϢH��1:k��t��̎��^��]"x�[Y�S��E���D��U�Cl�wm��u�U#.5�_H�ܽ�oU��i�)yI���(W��lƦU��Ky��0�.n��$�D��c��ݑ�5��D��9���)JVI�6�Y/g��Q;�g�l���-����W���խjww}������-��$x�϶a!�ې�>h���ߊF�a��TdM����}�Օ6n�>4졸����ȼ��9�8�j����^��7�S03���]��U���ͮU$���`c�<`�?~z��r㻘��6��XW�{i��V�|O�Ӓ�'ۿh� �*�[�L��=.�D��@�w�R�#��VJ����������ӿS�]�N1��E+&�f��͂��N�i�ٖ��m�8��%��E�Ců������_����؛-�v���YB�vZ}q���/rQ��>����q�@ާG��c
�S*ٛ����%�g�I����kn����Ţ4�$*�_��J����G�[6�F_�d���WٷwQ�W::Of��p�9��.���/s���gou�WEh�--����d�C��j������6p3$	�C1T	�u~)�k��\i�˳&�g���t�b�h	/)N��1pu�@r���F���0y���BC�����?��,�/U��ZZ��(KW��b�O�g�6I�:CƷ���{��1�aʑ+Z���]4���>D.�_����gD�谏�/�l0�'�x����G�A�#�xg7�{
�O�[Y{���M��[����#P"$ـ������a���o�uT5��vS���,68U��6��m��Ƞ{0�Yrj43 �]��,�^��rA��p#�k�;�����Kg�	¬pD\W�Gw@Ȯ��+Yk����0��.G�"�s���~���=�?�`�	R��k�
#�:DEv�(��G�~��/ə�ND��.��(4�ӓ[��U�m،��P@����j=<��ks��R��h@�VO����i�HDE�T-��;v����r��c�J�U�/�9��	+i=+ M���bYsv���k�zT�!�뙈vz�6��5ѭ��v��]_[4���W�jz�t!�G��T��k� Lۑ
��I���d ����zK@���g�LD4��n��
�6}�3��}�['"��v5j��Ug��_B�ڹ���D1�3u{.͓�^j+T-�/]�RV�Zd�웟�V�����c�L�c_�6s��ׯ�"۸�Hz��uU@����K�]������j�.�P]�'�V��N7�ga�<�O��ӒK�X�/3lg��5�±���*�cd��BVul�5�d�l
=�K�f�mzyr���L�
���ZZ��h�Rj.��nl8���҅g�+��.�ޝ����u[��.�gu�g�x�S�6]���ߩl���� �n�l�o�~="T���ùR�'��?�rú݄�Δ�o��!pm�'�����,���� 8�q�l���Qa���յ[�nȱރ�X��t)S�-�nbk7yKF�*�s=P��Q��z��4�h�����`��|����pd��(ӲD'��߯�m����D�x�����@����&>����P<��,�1F���3}�����Л"����#X�������'���JG�j̜я�K>^� \-\�=,������b��.8���3'�mt��8�{�ޘ.-'���uWƍJ�ˆĥV��md��@"k���h�u1��K��Ef������V��v�p�f|lRn x��5<�QW*��K'�@�@�ՙ���j��	1F:%�C9����wPt��{���R�,yW� ���͝w`d�<)w�LÊ���k�9�օ���ԩ�U����U�z(A�q4:X��1u?7	$����	r$�0�^��!��t�S'�)}���e�WZt�����O�5�CO.ѧD^U�KJ˯a���j���8c���cQ��u=��p@���J��w��S禊a����n��w�5�bu�]N6��ҁvs�Z�f�yt��`��X��:����vU���+6�|6CE�O�կ�v�y�Աn�5�g��S״L=h�Y�%5��c5�g�+0�߈�"f]vFz��V���̝:�4��6�^*���	��&�}Z��8o�����v!�f���S����^�'��؋�(��uB�����,݌WF�"�J� %L���Iv�h�v���Q���08�h�T��%^N������VW���"���9�2X�s|����f~:��+��e��/.(���Lɛ�Q��`N�x%�v,_�7qf~�����Cl��'���2l����I��)�+���ԩ"�D>$�h�i؝�]ĭ���t&M}²o�*v�Q^��\����׀����j
�>-PCp�<��������q������H�O:��l��x�X0]��y��a���m��=XH[��<�jtqW-]&EF���g��ATp�,/�݀n���3-Z���;��n4kZ�TP.�(��]����?��A��4k���Fk�o�<�"�3HC1�F� �a鄙��Q�(��[���}��,�5�	����Q����4��g��ͤ[yӑ�@�k;]�.��-�t?7��J��Zf�N>�jF)ƴ��}���~��<����Q���֬	"'��mѝ彩����²�P%�ən�G�,h��K����@"3���Mlq��i|,�/l�anj��@����E���VY�uW��:�J�̡4�S�S?�P���%��l[�g�k������ڴn�z%����/��N���o<��ɪ�[
��J�+ 8� ���-�Bm���QKwoծ��du����$���F������%�� `\�]�XkN	�ߩ$ ���G��}%޹�
凷S�}�Y����O?:ڵ�9V���N���X�>Md���f��2����s��hx�����E;���=�Oċ��^�^�g_���w-���H�g������uy�a"�K�t���BF2���Ҟs"S�p3^�\�ǁ��6$&'V2}�5��\�I&�+�YȊ\�E�]�:�d"���%m���>W��t�@�R�j�>Y^Ȏ��Jli�fw��K��=jS��K���;�Ư:쌑x���#^G_�8�Dt��3��#G�@D��>	�%1*�+�U?B_,�^.R�NvxгH����?%�r�{�I����3o=e�l�48ݵ����ۢ7��oĬ���aO��N%*���(z�R���Dm<d�4M)z��ۧ^�K�)7W�J��>f��c���kX���o�lRx߸/JV��g��Y���Z}�E��=a��-��:)�V
ɾ؏�j8��朒�l.���5����d�> �f�/]�o����q���&�|k�!�W�<�����ʷb�l8�P��u��W����
��1n|�J�韨���S�݆�`ś���>��u�}6�թ�xN��`��q6����w�|Z�%/��C�mۓ�W�?v�U=��鉜r�A~�Ø
��Z�bU@��ji���}I�`��6�q�/�0if�MlX�]��??���Q�6��<�h"��k�W�5\�b�o���-M�6��A[��׾�w�����*�Te���D����2+_NKw��VVzIQ�;-���
��9T�&aSi��K�rZlM��c ��XN���XF��e�Y����Rbb�����O����f�U]�)�)��:�'���T39ߑ+-O�v]��IB��2��u�h��.!����G�&�����q
լ#Ў��i��j�u��"�Զ��o�1qI��S�s]vX��4�g}�����q��K	���S�t�5�����������"U�L��ri��/�<�raq�{Y5f�d&�i� F���OL��Z5�-��
�7��VZ��нJ�V͇�	%*Zwqn���H'������	O�:g/7�d ��N�ݲ�����6{~���̫���8c�"Y\^O���]8������F_���g����E����^n��2nT̔��������j�I-+1K^�1���홿\O���RO���W��^��y��I��?$�3<���KΙY�n�ꗧl#B�XM�pKhUG��^�t�Q�����h�t���˕���n��as�-��#�`���i�C�ua`(�p
���C(�Ȱ�5�%n\x+  ��O�#gj\�Ej���K�Ԓ+	��M堥�~�`��e}�V��U�j�����䰿�y���OjT+���Eڱ3*p�/�tdӉc��$r)(��6 ގ@�4T_}ڽ�'��jў&��7�D��?ۦ]�j�m��%իh�-V%�������}�¿|D:ǟrgNƦ���z;��3��E"Ζ�q�/����0:К���TN�6�3���������>�u���!�{��F�L��n���`�� ����U����v-�5r� l46r�ؘK;z�b]4�*!�r``�(�1գ�i܄_n�U��U�i�}�0�4��/���r��I���ԗ���G|�h{�+=�M�b���E�*�Q4�y�{Ұvݪ���f�	���0ϵs0Zya���tu�q���&��qIC���T�($.������H��3N�_킊�*�v�g����Gu��\3�����Wx���J`���Τ��Q�֗+B���.wY��6���0�v�Y��S{�� (M%��n��Y��+���`�E=�$��e��Eö���Y��e����q�5�YUo��?��Y�l��8\�+�C��x�:2�}א���(�Z�?~Z�}ja�Y>��ϏJ��y�f�����5N�n��^��@$�_�	���:�T3P�(ċ𺫰}O��wk�����ᩩ��t��`Qgcfу@f��rm�bn}T�/�4%8��o��7�5�t-۹_}�JD��������O�M����v����]��u�V����w�(f=|9�|Fn��s�(��$�T���!�g}��+Q�^"�xܷo���k�m�%\�T�M��� ��8I��W�&��}U>E����+Fw�,�����5��';�@:�:q�m����Ł	��/�.�讕�Y4�(f-�1q��ƫ�}.�n��v�J���+�S��t��~$�!����Ŕ7-�qAF\��i����;vk]�8�879�V�/��.��q���zx�j�f���q�y�j�ԣ�t�G��3K����M�t��n�'P=Bf�A�[�}�Xm��(d���O�R�����S��P�	{H��(��x�����C�=1ګY�G$��fW��ɧ���!�$��w��FڅQ%��o�x��\���e�vp�>�r��s>TS�B���Q�3��I5�^7,TRL�|{u��m0�1�l{y��Z�y��?��dĬU���Ԯ>/u:�ɒ̔��^�j� �ퟌl��p1�^
x�ޝ����i�8.�=О���O���{5������0�ʼ��KALOEBOMq�""���*�b�,ed�m����G|o����j)slW�Nh���L��Oy������\���~��w��r��~M2SsU��;j���^K;�XZ������u�"����ޚ=�e��U��}�8�.���+;J���X�� \�^����[��kF���b���KB�k��q0�6�P}۵Y5�5��l�6��▱t-�eG��5�l���ژ}�\����}LҬ��V�E9&��m?)>}�(��Uƣ�;��b�'���gW�:�qՓn��/��!l\ܣ�3
�Y�����[���+x�Ys��;q�\g�Q��"��}��)Ib�Iqa��&Ȁ;�����H?��{C�Ϟ���Τ[�j��6-w�����V(����u>��� pE��ܞ���\ }���68s�p��8!��m1f�m��:[d�0�p��}ei��=m֩5�4?���v`6<:��j�^ߙ��	q���6�g��!a�@�p	{�O�Q|8�#*���	�U�����z�6h$�1�z��mC���������E��>�7����9�����G�Al���?m��G`��S���Ye௵Ƒ�Ы�m>�:�31Ia2�߳��w.?���ڥ�r��k�qqU_����{B|���(����j�8�K��1u�~o��o�W��3�w�	}f \iL��l� P�y���x7t�(�X�s�J�=j3��
�S�-ksg޷�4�A��p��-�0�ʎ*O( ���K�R��Y۝��j�F���3�dk&�Zt��t�ӣ������j%J0e�v��w���������U��s@��Y�z�6*@��=�z �ѳx� '$����z�k9-����M�TcA��52��h�"1�9y��6X�jQ��SG�"�E�!�_@��^C��u�_D+$bjͥv��^��M��i�1-�i���5
Yq�#�(�V�䁈�P��l���\�gVc�u��S9�%3hMf��
;d�d�UG�SM��x��<��1��Y)�eĬ0���G����S�5��[Ѓ�i��l���h��3���Q:�]�Q
>r��&shn�b���	Ki�"s�]�rx������[�0&�qxG���_���5�z8`�w�3`cU��g�ɫ���[�	2�X:k�.(c��s�ܔ��-�p��h��* ��+ҡaV�Xº��Q|�ފ���fr�eN1Fw%#~o�[����_��R�[�5�㆝�>�@�(pcd�G�(�3t�H�m���#@�u\����=���D�|D���dݪ�"#fl�b!��]_U���a!�Ƣ1Y^��a�)!��c+��:��p�c{mKne$\�B쳸��5���-b��mxJ
6��l县�*�A���|-R���Cycږ	�n�G9fC�s i}���#�$z��}�ad��c;R��QCr3.fq]�6tm�U;>��rt;�;�"�G@�?�,п���@�w!���c�X,e?���򉨛T�f�jN��T>�����V����?Ct�*.ʬ+k�����aU 8<Aِ?���İ�W�]�wl��5�����5� `��*̲�a#�s��<4o�x�s�d�Ѐ�엎�����M�}�`L��9Q�~ܕ��ePA7��*R��g��& �.�!G���?����]=������S˂7a�A��!�?�!�� "2:�De���C����J��P������{9~��ʣ�<ގ�@'�?Z3�Ya���X�ݶ���ڟքH��(m�&S���9���l�fLH,],��P�?����n�$WJ�ʑC��O��ח��;�<�A~~t@�Г��q�w�?N�
*�T���]��M�P�3Ф��E�E�_0�[���؁�=�������Æ��J6���)�%8Rt��:ݫȑ���|=���R��߽��x��ޟ�ͳQ]>���#�|�CnZ���H�c���aoy�6'�L���t<���!�F���T��.�aň�}�m3��v�t����}菺��ށK�Vo������hZj�\������|��a����� ��D�4iaE�v�f�ĘD�����+�!�Y��: �V(�kb�4�����XA�b��_��L�K'ܐZ�wF�����H�ʿ�*�r�4�hl��M�_yÿ���v�g��SZ���e%;MNe !��A�x�q�:�4���׌\���[e�&�@��I�4�VC�lK��a=3�.�7�E�N&.�E**|ˑ��`[���o��T�\��s���;o�Z-0�(���&s�\�H�ge$�+�f��@@�$&��g��U5�f�A��e�1���;1�6ĿO�� �ޡ�+����ˋ�XX�Yl���u��:�E"q���0�R�-����m�b�ӫ��}l�!�����g�ܚj*T��HUz�N ���~������Փ�ak5:x���y�I�ߠ@i�Af�.6r>}�w��l,���'�h��}c8��K��ܵ����i���]�oq�3+/Md�$��}�[||��,��.���u�S}�b�Ȫ���g� Z>����m�;������z���n)�w��V�]��t^Wut�O9Qs����N��s����C`�=����CD�����Y�#��Fk�Q>#8���������N&���S�J�/<��fr�g�?��l'�c������m�$���_�sٳ|����8����f4�ʼ���V��G����W����5���;B��{2�L�t���������e��\*�2Z� ֔M�"�)Y�?����$jv�F6����3�Z�p5'��}V�'��*�(dd��� �+y�JG��E�:���;DR[�%�@��n@��kc�����r����A.��1XZ�d;��f��O�^6��xM<��D����xlG�e5h��R�E����*�A�h�'}צ�`z�-�%��H�m�*��u�(W�v�ddzC%�wq�9*���V"�̭N�c�}��*�gxU�.<z.��^>g��	J(5Ѽ�ǉ��H�YNY�Y�XT��h���D���"�k�+��8� ����F="�ڋ�1t|q�Y����a,�5㸟E+�u>�3r=A;���"���l����|	Ød�ёƫ'�_����d5�F��g�<J��+ϗ�`r�?؟ECB#�u]k�d�,lbpt�k�އl��첄�ʘ���p�Lz�[�~ؼ�p�?�w'GLϊ�]��e�b��+�\1K"�^�:B&���{�>� �PRS�2�0��**����<v&YG{Sŭ,��cr�P.5�qW�E�c2(z P����NuGܗE��@<�3�4K�߱��1������߹)Y_���[�c��V��RY��̞9[�Y��H��m��X�¾���=�mV�gs:��cԛ��5�����'�iÔ����(WNz�����]!�s����6�{r��ߙ����d �,#������
7��#��;*u�z�GC��HE�U5�8+�awf�`�y��i*��nT��ǡ�~��O�����E��>��V �'��6�L���Å����W��0����xZE(#jd��lf�פ���M{�����P��>n�#-��X+V���Y����1�����(|����?��o����L�'ƨ�b���"��II}6y���EM	��&�k��_	7���"� �l7{P4gA��xw{{5?���&�]�^�#��nG���G�͠q����3*puxݳj�H�<�7���O��12Z4� ���i�Kzt�6�
_6N�h�z���9t#Ȫ*�� �
f�Pڭ
�PZ;�E��
)��l�!|B}@U�F]�w��J;��c������{��aBj��$�(�2�V]����{�FW�l�G����ʧ	��a+߳?h����+��g_��<�����7���GO��.��f �H�þ:]d��1��x�gc��5�R�Y�^�v4L��O�,�l�д8隗3�E|_'m\���[�7n�}Y�u"�J<;60�B9y��jß��v�A}L`�Й�E+��_ڶ �]g�H�����Na���������s�WR%1�A͎�h#��x ��V.Z"^"�X��v�*�a��P��S��S�9�> i�۔����>"U>����ᓣ���=_EW��Q����פ��,�sC@�O=�]������:�X%�f@�V�7���.<���'PU���)uIJ���ŭ)V���g�`V���	�d[��ˎ��"��O���&�r�6.��E�dP �s��h��ֲ�:������h`&�Aѯp�yd|&C9T�w�M ]~�c97\����g�n58�������)�z��w���B�қ*<?�yn�&
�]�wQ�#�ƴ�i&��u��^�ezѵ�5?�V��u3ࣶ����޶O�.�a��g-꼅����:Ì�߻�Ρ�ye$9�ށ�> ;j���`S�4��s�w74ˈ��"+7�(�ny1z)�	7�h�d���S�7f��|��z�k��l4���? 2:�?�&��4N���ox^�N?�ͤ�q�8cd,+fD\��;'vA+y�Ť��/N�{k�p:@G�ס- ��t�U+����]�y����x8��Ø.����`�|]�J�Y�~gNR@iW�J�Sv]GeĈܙAܨ0{��i���f��y|Є�@�ޑĤ��T�1e�E�6�U�T���H?~�ȴ�r@P�(��>*0����o��y��〼��m�r���A|���@�eu��kY��`4_����D>�aJ0�}wc�!�����q�I*@�Zz�mꏠ�`��4������$����N�rS�H��޺n�o�O�ܿ�.f����,�������@�l�K�5y��}��~�* WЄ2�~�~6��I� �������Z
P2G��(Q��7>���J�PA�����OGn�*�������Xej�������Mp[�>h�[�L�E�-�_���f[�S�
��E���?��)�7{B�6��0U�n ��;X�2�5N�<�M馓W7$��  �NC���B)��b����k����7]1���X0�߉%�`���ߓ����D��1`�r
�4�:W��?�w����G\��{o�~ ���F%Y?��H�<{�ccW@�� �W���8,:����$/�p5p����le̦zx_g��{x3����CV`� Z�πx'����f@�BZ���_�c�B���݉4f�[����@�����,��O�>"�����?P r��{����/���-�w�<���9���AAq�	�Y�[���sO8��M�!W�~� ���c|t���xFm��LɊ�2����{n(�Pޣ�<�Q�H2
�H��}���y����jϞ|��u��s��WD�{�*�C�Y�D�B����X�<���tS]���ׯ���s��M�����O��y������Gm�l-�Q1H�e�_���K�TB��E\��D*%�Z�l}�w�"���8���ȯ�Ro opt�y�箣?�{{T���E��,�r��-T|��Ro��1�is�V�yK59���n�n���B�r�Y��? ��.i1Hj�'�]��g�f/p)�PT^|���:��wlF�Km�w��w�$�b��P�9�ȕը�AXo婎E���C�@G����=�D���T���w��/!�T,����ӕ2a�L�w�����I�;i�P)Uݽ�{��(�|��̷yRP���"~�с�`��2�%/����Z�XVD³[|;�� Es+���)? �Z/C��q�'oo��X-�a�4 �n��I��`�	����BXP>#؈�9rZ�R+���w-I��D�^p!]���#��J ' '�ga7��܈��'<Ac���|�͑�UF��-��w�b��4��.v,�Z.�X���0z�g +n��g�3~;G�I�v�^!��F�2�$�.f��0�*I����"f:�:xU�'T�8@3J ڤT!���J�P�v=P���������	u��p�\F������i�:�A>�ug=a��]z�V��?7���Ř���BxR��g�YInA��I��a��)rL����s�]�Vh�$�t% nD�w#�;(��a�������t�$%��T|�խ��Wjl-�G��g�PM�_��ڥ���-����NoJ3r�j���S�冦ş�\#e��:�Z�ny�so�J_*�Z�,���t
����ߪ��T�Ya%E����T;u�s�B��׷�qq�����
�]Pu��߼�?��?��9�0,8��M�r�쩕�g��߄I�x��9 ?u+�w�S�G@E�,S� ��|JG�	�#�i��f�3-odY=��c�R�0������zӷ/��-é��щ�����G�<]�1�SC�P
U�;\lv����V�
Hb�O���<С��P=�5Q��P��@�bi�xW=���<�U������*�:��~���VZ�gb��F���Z�Ã�V�AFIO��iD_�a^y��$��Ն(/;���H�ar��ۢ�󳝡�-Q������{��Q�1@	q7�1�[O�\TN���%��n����W���I�i��j���G��Z�;�������\� Ϧ�THd��W��WD�Wr����W�p�����ԱaG��+� �vP��e�z����tK�]��Oh!w��s<t�Y�z� $��R��1`K�[�-!<N�"���׮s��r��N����@���*�Z�Ƹ���;�Jr��R�Y��".����{�] G�)�Y�&�3�ݣ��\���y�I���l�j;X�K�_`АǏZ7��S���%ɪ@|ו&Y}����T-�>�*����#��t��jԄ�2(��<h�pj�j~ew�<�X��N�Ը{��A�?���N������rzs�\��]�.ݽŮ��� ��ĎY�@ދ���=d�dV�DB�w"E�x�;��b�m�>��Ȕ�wk�����\<\V������e�8��+9ۀ�]1 �>`.5Bvc�yz��t��(����� �/�oB=׬��K�z�DH���!-��d e����H�q��KK�^nw�8(8�D jM��MU����UKݴZf���}GCY��oDmq�F�+諚�">��$E5@猞�̇:���V T&�s&1 ��2��Ͻr �;�wd�o�<��x��{�t�[ؙw���)�Cc�?jƣG�q����q����1�K"(1ea��?g��\�Q����e�3��_�e{]��''�j;�޺�r�3��^a�o�$׋��A�L'�������@��j��M�	�&f=�g��A�2��c�21��<f�,�݊G��_�R��evå���5��<`�� �b��]�u��[�E��$�Ý��48j�ӌˇ	ر��x�&a��2��?fղQ��� d.M��tE���*��#��>ޅ�Z�\�3p��cVՀ�o�� �	���X�Do����i�W�,+&̮toڹ�f���hC��8�dBT�D���UbP���t;Hέ%́l)"V;���NTH#�`qHgݼXT�P�9b�L��Ru�3�&�-X�*���R��|W y�fG6��A����vD�.��wa�#"o���P��`�G�Eq���\7^q(�2�l:�m�"H��S�[��g��u�;�񅽉�� �,���t��D�E����tMrk����q��F J�_��p�8Q���L�@��L�(�k=�X�4ÐA�aҡ�#����{��"[8aQ*�?��^�k�p�r
?��ަ�71T����O�o{�+AJL�hMUz��zh��`Hx���XT�;W�.JH	�2���>RR�Y6)2����b�8�
X6��(k]V:�˴١������J����˰�����E�FI#�nmӰ{��93�1��M�"��K��:v1��Y�j4R
U3�X���jى:�gN?�뾞s��Obe�SH�M`3���k��JR\�_`����d_o����GF�a #OV�K	�'�	������_7`�. ��E��@^z����:��c]rx�K��,����P
��?J]��a2Gw= ��kY�{B\/L9'����Ï�OaNx�Ն��Ʉ׻�Wl[�@�d���H���IS��k��ٕ��/B_Q½�J:�N�a(����+��fR�\��Q��� ����Շ.�@�����)�i�Y)`�'U6Z��OX�	�J�*Oj:�a���ɧ �<��.|	�1���>rPT��
�#4s7C2�H���7����b��%�V��ّ��}�z �����J }��L)dC��9m�br>
FF�N���[����?��L<�%��t�O?���@�{`i���� ����Z��2ɾF�w8�ֿzv�-dpWJe���!���^���q�q��c�Z�6�ڀ�%�JΎ�LA����dRO��Iry���&�ѭ���Q���r���ddAd�畡����0W��4�y��k:�Ķ�Y��r"�n*��C䅵�Ha�¦�C��7��Fo�<���N���9����,} ~v�I�[�f2���Yu^�����wö�J\t� o��4��R��o. m����P�w��_b��3�n��tH��ݡ���?���Fn��\��sN��8���C�v�%��������凿�����Ѣ��Hb�ݏ����LE�'���պenn-]x����/(dO�}C��e��X�O�Z[�4��@�#�Âm�T�y�Z[l�vcn�	���؇$c^du,V[�{��2ΐ��{$Ve�3&p�l�ǥ���3�� ?�۰ԃ�3.\��օ+�(���:O��,:��,e�������-^e��Zk��-��k�]�<K���i�S3�s6�|!����%�Ǿ��K�Q�-�~��4�0�Wzg�Ik��I���aZ��g2γw��R@�ĮA,������;Cw���q�\���?n��%�C�}�y��X!t�٥x�Q�SN�j��*o��D��]g��r�8ӭ�oH+f�+�
.<;d��{12?��0\m܌���]�(֏�V̗x@���?@0��,ծm�5�,�Qs��'e"�0>u���Kf.�P����\7�J;:dHk��7l%��"y|�ݩܿ��ي��l�,��Ud ��7��{�+��	'?�1��Lsi���",W[�FX^w�s��v�ƺ�嶺�,�n7��Qx:Q5c������0��[��P1� N�Y�o$4��n�yd���2��=�rm�� �S{!!>�L�$�Y��}�l��������]�aq��!�I�R��>����Z|�o�W�Xﴂ3���SSC��e�֗�]��9�D|��f���ʧ�Q󹴥,ΗS��x	r>�z����=���3��E5k�?�d�f՜�~�a'�o�H[l���9Dr���4=��*��x g���t�M����j?�z1�:���)���|�5��}}.?�����FZ(�K7�O1t��2�?��'`������O�����h˘�T%�Z� �e�ϖ���:���I��D9�,�-��'>R�G��Br�����#��X�Dh6RDp���RF^@���M�Y��CO����߼�j,]E��@�)*,���*��0���S�z�1`@ح����{ǆP쾩c C��t�ܝx�%T��<֭+]�0��7qz�q}>�+S	��\��ю�z��q�1?R��1|L��P�cK��W`0��H{?n5���`�"S3W^"��")~���UO����n;�m-C�W6��e��-�3=�p46�޿1��/��xz{հ]<�w��3�@^gY�nh�۔��ME���۬�eex��;s�>R��Uc2�c|�#��L�3�_D�n�
>����Wݵ�9�x�+�'����9��#]MC8�����\�<wq�I�|Lc�b@D�p��v�W��B�,¶��ǯ�6~e/��O=w͆��1�� L��k	��&�hS����Tyk���~)G/S8*�R3���a� 	�R-�^.�� �#�0G����Q�0���ٞ�y99�Hd��-��]���^��r��n����HV�	��B��Fy�Y��G�8͎,���q���e�k�J(A��^�_�L�uv�X]�
���@P���Knd�F+ڑ��(՞Y�W��68W�!�\�H�������,����������5�隓um� �<q[���C��d�,@M�} �S]���u��l]x��^jJJ�g��4�W�����{�mq�	���;�����I[c�T�_T� b	G��`�b2�i"p��O�E�k$��!7ʍ��
u3εRǸ$�|��:�`O�`i�SK�E,{~2�)�+C���٪v�m����l�n��Nf�C�����g�������}��fz�P ���|�1��+D��G�S�un&�~����5-#P��E�\�m
 `��;~<b]�����t5������]K����"�<�&Fc����
�郷;b)L�$D�uE[I���������I�Ӆ�7���e��3E�`�K�H9�ۅ+�z����n�y��:\�mOس�^��'H�ޅ��G7�_��&�6`P�/_��J+/�Su��M��M���;�݄J��py�����^�l�9`���F�}��[��/��Ӱ�5�YG!�W	3��nB�}�L�י�ȭ�$e�֣S��BZB�=��~�
�̥�C̍kn��G?f�Y���zt�����`��5��J!��\����Eu^�����0�TE���<&Q��!r�M)�����]azS���N�;��"��H����`�\77�#�r���3Fq�<���*ЎE7���_LŌ #�Ǹ&Wy�W�QȳԘӀ�)}[�W<�ӟ��Pm�~=JWn�$�27��+��ȳ�$7�U����N�$A]r�CSBF�&w ���T�O[Q���E��=��=�#a��NRN����B��I��8O�P���l������
c�1x�t�~jR��/�oB�c��s�҈�4�����۰p����S��l�P�h��]��s� ������6�>��O��k��y� ᫘����_q8���')?J2�|i������}%̺?n1q����f�}��K�������7�Pڗ8R��m��+_�D�b��}IFp���}��Xe�/Q�?⎙��-��X��1W��E 5��_o�vi 	~Bk���7�#�X{�RV�S����7|.z3Z^��%���~k��\���G�`�&ːPc��LA_E躂G}��b�d��Pγ���Z��g+Za�D��$LҤ�3F#�}����fܒT�����K�cc+�������q	&�����2gyC��B	&�I�g��|z#7-��;�+���l�Jy'�P��x���1-z��������I=�[]��c���3V�Z���452��k��{'C`��S_��E;���t"�(��2�t���t��HJH3t�Hw�Hww	C�t�{��{��2g��g�Zk�{fƜ`j���k�9�)�稴�fC <��{��I)h��f�g��Y�=�!g�,F�t _�6��pko��$X���b,=z"����ԯnf��R�<_�yM�<�a���z��bT�~��2Z^�h�twS�E`R	���T�����r��${6bŇ��Z�i�S[jR@(s�8G�+??�2!�7W��֋��/$��ކ��ߖ�GoP��� ֊�+wc]�i�.��5���q&�b�e_��d��"'�i7��:B �-��H�@�P�_0t�0 �J�����	�s�lwu�6<>����v~��8M�{��'J]Y�.��_�Kw#�C�?�oai9�U9����"4^");��ݝ�~�b'UN��	�ĕ��<��)�m��0X����$H{u�\��������
d��Bw�QF�6��V��>�Rw����Y�\a����=��l�ͤE!��Wn��ڵ�`�1#��k�1�y��cP����&�����Fy��n_�����4HKF ��VC=�K�np>L���j9�ȩ"5�C/�6Ө����0��Ð��p&�f�S*!�ک���Њ��ϖzE������E Mv\��MĴk����+t����$����]��7ֆ�S�U�9��c�6��xG��|'\Ѝ*=(�u{'C`�Uk��~Q;���=�t?���D�x�ǻ�T<�{ƭ{S�5�1��ce����D��|n�k�rQ��Qn����/	�`E!`ŔV#Λ R�@����v�����O5���P�p���Ȅ@\���V�7���o�YJV���I����l��8Ј�\f.�Q%�6|����u	{�Gn�n�r����g~
u����呥���f���M��1)ۂ���o�V#��W�0����ߢ�}��^�L+t��54��/��xA",ŗ������f��o�+�<��^}�W������2 ��|}�e��L���l�Kh#&�7����6�����O\G�#d�'`�ԋ��ZG�G�&+X�����8��;�M�.`E��A.q[�&�Oj��E�[Nw��^%,��j(A��-&�,��,P�j���83T��4��C9y<u�'�C�'.�$�XM�����g�2�|�N��Ab�Ƶ:7Tmł�$��dy�u�˒�L���<?�o�K��ƭw~�	�O`G|Ά��g+k�k��ۚ��E��/��쬔��s��CYڣ�E�_����a����nS��Ae��2���	b�6�n0��-k�r��HT�bɤ����aθ�j�%BI�Zp����C�:��(��~��T���뼏Y��@��
��,��pqk���� 3	�r�������D9�{fʴ�#�Z�K'yU�h7�_�hR���k�H��_s��ǜ,�+��k>�B��~��A/��ԩ)�$>t�,YxK���}�z?��E�ӃIinp%�J�c��{�t�G.��kcy��3e�A�|�!��� J,�կ+ތ�Q=�`W��@:�z����y���\�]�9�~N���m�ڪ�N�*OEA3�Y��;��o#���H�S�|׀ד\������-T�4;�Ş�`~��e��FZXN&���Z���%'�S���+l�g���=����t�<��G]�B�dA
��/��>�h��4Acz��Nr~��=�g||u�^��g��?`��P���������#��i��x����qCU��U0r�\��U���tq��xəf���^btH@�u{�t"�%��5��?9����<��fW�l��R�����7dT���+!ұ?�%���>� ��j��0]�ei���أ%��r&�|�Fք��H�mO�� ٹ��w���?�]�&����$Oa@	J��O��r\2V�X:&��(�����i�5��K犯7ʍ�Q��D�
k�k�z�k�_Y��kW�%����r�aap���'jȈ�Y�噁���<oW�H��7�nk���b�=t�S�h��Q]�����VE�t�V�Y�s	y�P.�t��q����@�Oy�'�b�V��o87=�'3\�
�5�'���[�u��M|O�uV���|r�Өx�}y�C����g��ڐt��!��cŞi[����9�ᴯ�k�`�rS��I<',/�d6��6WP:3����Jz1W	��`p�L�v^XX��SN�V�)�!�&�f[��ezC�T���3'�`6%)����^�eQ��	']q���X�Ǥ��O�Yu`qsT�����\�12&�=?^�i`�QW��=��3�C^��Wi/��QbKmϞ�S�n~�g�s��=>���?t.A�CiX8�t��Y�h�|���n�����ᓸk�{����H��O}Լ�{j�GU;O����-�30���g�gW����^�N�"3#hW�|�~�
�H�Z��s����(]��{��ǖKY[+�Su�p3F��<��A@�����=��3�����D�t5N��b��6�Nc�~�d�N���h��g��u�����}r��xNJ���v=j{0���7�u|���D���P��q�.|}�j�L9�������
�_�jb�'F�$W������oŞƩ�q��mw�� ��.���8�����]�Ac�eT����	��Z��GSl�s�r��%������lug[�Z�N�����%l���I����gb���h%�n���D�=��y.~��W��<��#=��#!��q��&��n{�l �_S���1O����]򬞚���O/5���[��o�*�V!Y�E�x���%�=��o-;�6�VD �=��n��œ�fH�&����z�$_��Fosf��ص��I\j�4*�C��������\���E��&)� ��bvCds�zj)��WD�k	^I~���ye7�
�:ś�[ݎk�H��%��Q�^8c��� 3������5V�'b��9`,���#��3��[ޤ�5���҃ˏ�/N�g���U��kE��b�F��)�e�D�$y+,8QVo/�~�a��ۀ����E��Gz(��{�B��"('A�����^����d#���R�g�j��D�"�i/����V�9�4����D5,�o�< �|��F�� �!��H/�aO#�&$QiMe���*;�&C����a�oJ�	]��K����q�^��2�B7E������J���Q(����y76��3����y2�f�\ ���#�V�Y�]9zN��g#�k��06&g�z~Q�o���P1ٸ߆��Q��}	�:�wQ���1&���(���$������}I����K�X��KFQ���W[b�O�볯��?���F��<&a�喞�]"U�a�I�&�L��`	�$�=�Y|jڪ�|D�������{�zǳJGT3�'� Ւi;V�ƚ�X�� )��9���<�z���2���9��a9���#�C�5m8�35R?d���1���j8�ga�!QP��Ѵ�!&tk:�*���8�al���n��I��~�9<����mq����վ�ϵ\�z�C�8�HH�s�`�E!m�mB�����1�����@cT+	�O���30 ô�q��P�Ȫ��ﲥ�&}CN����|2D��l�?M�]n���h��k�2@Ȣ�W������rm{O ٚ�0�'/���R0��*8�3��WE�m�zJ������7EX�?7��g{���ҙ}��4����%Xu]Sy��ԡ��P��`0�9�_~��}&֟#OS��>��񸯤�{��ዶy^ZE�D�1z���e�>v�E�P9�
y��xg�ys|1+nw;����^$����7�}7��2��0�������Ͽ
W��Hٺfi�E�9���Y��2.�}5Y�T��־�P�y�����>�;������o��;o�G���i@"��3�Pl�1�9>���Ԉ�ܮ��3�b�,�>?����ҟͨ[h	�v��0ۏ��HR����He���檌l*O7:��]�R�u?�9�} ��r8�tչ�d�~��x]��Wө�x%�-_m)�|�C�����9�$m�Q^Pa�*���%�����I������qɣ͊Co�³����]����p[����D����|��$$�ҭV�|������w%���:c�25/��@<ёF=�:��j�c:#�Q0�����a��H��_-����!�ji�-�j'����?�����d�wݥ�������l;�j��[��oa�˼����:�Il���d_%in9y8J����Js����9ʠG��pX*�s���y�!���IL
��}�4�r#_@kh�L�����V��$_B��+���62���t��n���������2��l!���bx�I�z�H��n�_���M���/�)��*��Bٓ��渼�ʯi��J{{�[�[��r���M��n��?bO��A����VA.�"��wy��g�d������{�HYf����a��U˧�ǒ.VJ���~G�4�w����G�ڏU?��{bv0k}%ګ��#
	����(/�r�]�_)�?�,��>���ϣEdf<�қ���0es!����U�.�M�Q�)��]^9k�b��L�6X�zU4�r�� ���?[��X�|k��2w��ɟ���~�IC.�#��7v���Jq�WvT悥�
�घC��
�'kT�-Ё����E���,�ݓx�gg�t������Y���i��oB��efi  �����蹬t���R�-+��NՏ#�
s����=����ܸ�;P6d��YNVrhĈPI���pO���Kvc�Ȥ�UX&�w@_s����p�{^ׁ�H�H2N����C��ēƔb�z.��f��F�N��z�\n�'�CJ���3��s��ݭ�����Lv�Ή�h��q��y	���=l��K+AKn��2!p���jn�� �@Dx]�d}_Y-u��m��2��Z��Qǵ멟��eM v˩�����*��͉���(v�y �6��Zf� �r+��:wk�+��
B������t��%�U����Ђȹe�W�C x�'k3�kXJ
D�ii 7�%@eg���ʥ�
�!n�;�0\��!�$OF������{��N�7/�ޫ���A�H�3`٩�BG��M�����
&9���l��ZG�	hlm1z|����/Un�Ԯ�Y��ݝ߸�p�8Q/P"jg2픛�5���f63��:��7-�n����B.�k�9�\�u�d77�8coz�[뚨hWC�VU1Ӎ�bdv���U����WTHFw]#�`�/�����N�ߤe3���>[;L��ai�R�?�����������ۣ^&�琗��笫�DT��=Y��2jz�&N���H3i�=�'M�.q�����$�$Q����:;w�&ߴT��j�kM��Kz�Ǹ5"a�ܬ@94"pg׳������OK���wA��5�B�x�rX7J ���!g����&A���I�i���|�{M�a��\��H�Z�<gd8����ϻ4 �w�J���-�߾[�P%�@H�ۈQ䘶�GD��v������D�����e2��3������Y%H�)%��a0�yTwr&S�76 \z<���
U����xt4���O��C7Bؠ6w�Z��?���[ֱkw�{�G�����o+׆��뀠�������!���/�C`}:, �v*��Έ���D���h>�c]Nt��(H��,�ͰO���Ԙ�ID�n.4��՟��[��C<[}P�^���ӈ�� �:��+m>!q��$�v�U��C��#���si�?�����o<�ˢ���)��\�/t�ux�f}��ֹ{�I�@�Q!'Hj�F�
[��M�>�q��/Ƚ!-Y��[���]�o�z���,���aj��QȻ��m���|;c_���@R����/ϟ甐��4 ��F0��À��,��p�/{S�L��8X$�?u�~����5CQNN˨ڴ�p5�bx�3�='����K�Xx$�0N�G[9��¬S"��~�\+�<�R�c�x��; �>�(`��66��9ڱ(���'S>�q4Oc��eN�,�f�w.�gy������z�6���~#9��Bɬ12�Mͦ���*]%�E��h�;E{A����cBnɻ6�fGϰ*Q	i �F[�?=�8F�-�	;���]�_��h������n���I�O���Pp���ogT+�~�����ݺ�e
�L�^M!�.�"���)��5��q-�qG��$��hL���<�A�H���3�a֨�R�>\����3����nz��,��E��,#�^t�=u�, �!T��m#F���@f�]�;��*pd�F2s�{�x��"�2Zf�g����Q�|�v���IuN{y�Ϙ'�Ȟ��?M ۑO�5C������2^�aJ*��vߠ�Jh*[�P��Y���������A�#�k�t�ce��2�R�� ވ�;���� HUx8Gwq�]���W׋�vL��9��NU�T�f/l�u��u����Ң�jG�]���KG�-e��r�?F��;�5���W���B��5X����[��b�x��?r�l��kG��䦖���çi��74�0�U��C�\�?�F�h�k&b^���S
 � ]�Ǹo���~r��@������ D��׮��5��t=�洘��Y{c�U�b	�apnmE>�F�c"�}M�Z2�WU]鑫�*$ �A ~w�X���ujr������j� w
�|�֠~{�m�H٠�<o�h>�g���Ex��j|(ݖp�]��4�������ϸ�Y�1n�}�T�)]k��Z(-!�@LmR��~f�/oHٗ;�B�&NϹ��U(^���xY���kV��Eer��X���� f�m��xAz��e�AW��W`��Ů�́ـ����c/�2�Й�>1��K�z2�6� �D�uj�sg�n1�o�%6��8��ZWo��̏�*��'
�>��͊�RՀPwT/ZOF��8�,�|��@��Xh��6�K���CR�#���h�[sdFĻg� ��(���^4�� p�z��z���8�R۵7?�!ꯡV���@@�n>/�!!�O������И�C�K���[K��<�3�"�TOc>�����iql	m�oo=�j����|��pė{@W T?�����A��� /<a�	Xp�G�d���X�E-�"b��G�䂊
��:�����~w%�q7����6���"v�~�,Jr�j}�#���;L�V��q��2��q���Q߽Kb����i{�Q��@4u�z�����'��'*���ATYy�vp�M �*��e�,��H0QZ�Xu�!Bg?�@R���2�X6\�(/��k����B,�j1R�N�$7o?j:���Wxq�&F`�7�y՜��]��Fy!�2�ڃ���@��y�oot�_��?( �������yt�F����3�6�4��f�O�����A�h��,���:Vj@�A���Y�f��Ϭ���y����l�h4���uX��s�����n1[-�jA�l�"�r �rwG�I@��I$r^����&ށ���~���EJ��Aa-9�ÄV*]7�q:�}��N��v4(G!P9�B6n;������x�mzȪiIp7��Z~�OT)ڜ�3�uʔ�6<s�w<g�:���x�"n��0����7��u����-5Ek�d��]���ˣӌn��h��Ϥ-,(iSt����%��������ap�˻��el�2o�����@��it�/��w3<��F9!
���%��n��@a@�:@���R����R�<�yڀ�k�\:3��@k�<̰��A�����rǤ�374��~q��z��8e�"�F�vG��݇0P�~��
�$��THI�S��"8���4F�� ��rk6�I�v�S�ӨC�j`��/P������nO����$rs�p�>?(��%�:�w��6�8P����/��L}�;�#I�L�w��L؞���<�D��i����|�T�,�ż�M�nh�g\"y�4�b�G�%F!"��g���\��	�/,����6Sx��\c����`3,Z�َ҅�iTl�#7BT3�q�DUm��Y+
	�bF��U�0�0�5((t���w�`x�p/KG`�����S�W�-��/��YG'���L�������^y@���fk�".Nw���{З�j}ܺ41�Y}4����㍫������x��V�����8�~[T���d��o�f�cB��ܲ�}���-c	�b�ka%?4�������󭍏�і��@�l>R��&��t)ǯOh�!�&���2�0�� �N�������`:��?���p;��0�0;�����Z���u�?�_�BL0���f�v�_���OM��\%$ȳ�S�zQj�<�sA�ę���ֵ3���|�r�1,��@%���'\��6ʟT����?m���3��ښ,ѷb�q��^�AǎARmv�_L�O�ne���nn�B䚍����C��q�= ��#ϔ�6��������C1c�F�R�	R1����e%G�V�H�)���GSd�h�5�3H�n�|z�5�kC���E��C�='����h�v�w�K�r�o��)0c���"�ΰ�T�|���`(����\2�%�vڍˮ/���W@�L�?�|�h>9����:��ׇ�]�G%����.��x�6_�H�����Y��&b�Ƴ�@��)*i�T���j
鑈�O���<}Y�>[X uL�<�Hr�o�|�i��|LƢyO+��ɜ�]:f���^����kGwzY��_�I|( �۶�w��j@���їvRc<�l�ltk�)_���t'7��.9�;������^ߛ}����+;�zP5�LJ ����>|b��R�h��,��v��4r#t�a%Q���� �X�qGڼ~��Yj���DR��i+�41�MQ�t��٨#ԕ��>jO�Yw�#I.Pg�u%*����{����L�ȈQ!�و�����;j�ӌ9���8Dߚ�,��j�BҖ�ܺv+X �B�1_Z}�[vvs"&:J�h�����r/RQK���UNA�3 ;Z���o��lL쉏eJ2^�zO=�,�5�{j���%����� N�����O�4��{�&�؋��q�@l�#/���DNw����>��%�T�=�u��g�6N�4��f B1��"Gv���*	�瀣A�Ayj�� M&g!�;{Φ��i�F9���������|������X�f�z%�2�(<( pʌL�pt����w�*��H?{��V�=�5V@z!t�Kz�]�a$���1�[x�v�q�w��EA��AH$�=��B����N�s�)��(-^��;���^�_ qG;��a�𭨤i���[?�^`�D�a~mW�o���9�c#W����P��7�f���E5�ʍm��{��P>�xg/�ӂ?+?���%��T�|q4v�������]�x��.crܙz��5Y����sUG+:M�k7�����5�x��ʯ��:���	���ܕ���ԣ���� u,-S������V���6�C%��&��@"�-�X�[��'z���O�`�$7�:{1��zNRAΪٷ�&��Iy��]AoX��d0=�ϩ&2�p�EVU��u��Kнy7f9�vU�g{��ƑJ�,�����:��N~*d�<N�RW���{���~A�o�ΐ��y9��Y�UCE�ج���a{	�c`��x�F��?F\#�@Jޗ���X�)o��v���L����'�q���u���>�n�N���)^��q�TAYh.��l2�Iz)
Q�${n_Tv�Q��+�ϊ)��y~���Q��$v�.�uȾ����%Ewy��/�a)> ��լ�l��z(��oTb℁��1� ����qT-�����Hv�%W %d�zg�2����bV��x�Ǜ�O��ú�NR��h�<�[p%Um�
#��h'P��'������l?�GP(x�i�A�T[F�	�*����u_C�D:E���ߏ�Ph�y+0�q����ְl�o�!������V���s���M6ӛ���[��ꋣ=��^#��3�$�F�s_�����x�5<��z$�I�P���8CG��n��s��9���TLX�.�硁�'L6��eN~#���u�	�91��-�.���\0Ӷ_ǥ���x�9�ůhH��<�A����m�H��p�8:B��p�hۣ�=��^o
�⿸���[���.x�-�Qq7�K���r����3��Ѩ�S��zz��.3>t�/eZ�u�م��خLI@���p!�F��6�Z���K4Odx O=���t���=�<`�|O����1�ln�	��U� d/���a�D.�A���^)�D���ɰ�����9��Gdi�#���}g�ʼ��9΁ȹ� ��	K79�u�R0}�D�2h���X�H,�Z��a ���A�3PzR�&��v�y�G�y��mEM�z�q�zLpX=�~���ћT��}B� ��+�<]u��}5������8�i���{�g��Y�k{�����)2~�摶5�� �H$�:�)!�ҝ�S�ed���=
��x�J����"O3K�D3;v�M�� ;�ϳ�^0\:48��LvV�c���$������[۫�GW���[ �/����B�]��~E�SZ��t1	�稟�m�﬜����̛q47����oZ����5���y�f1}2p�������j��a�T�(��)?�E�oԢۤ�3<R[zK'lID6�CI��
F�$���%,Ny�~xT�[��&�6MRV��N�H��i\~W�3��~�'��� I��8񇔔Ժ�_MH���9�]��� :%%'��2_�Z���)�a|Lֺx6�h�->�,X3^�߲*
=S���ix]����a�ZI�CP�i^n����?�����3>��c�H����N�c})X7�+d��6�	���Z{�9��%�����\�(��JG42Q|w�aJ=����`ũ�B�ˣ���Fv����+��	�W3���G��ОQk�W��R޾7��h4ߕ�xf�m\C!�m���-��|�YuP%�V�0|/Z�����O��U��^8��d�����3jb���ڇe�p9�c���n	����D+�C�lF�|����&W����f�J�=o���4���z	D�)�VZ]t�C���-��;uƮ���;q �^}�2m9J܊���>Y��9� �A[�a*�H6@š2��V)�(4�zr2u_�1�����x>j��y��}�t��ʣ����u�9�1���A��o�X�|9~��1�'���fQ�P�Q�z<z�O�P���YWz=�/;A��z�/�<�hi��I�1W�y�:�w�Ŀ�o����ٽ��LoԚuj�t�_Wy��ئg[��X�6�<C�D� ����l��*I�� 'a��ʝS�v��/���P *ވ*����.��o����;�D�1D��_���늗�+Ƴ�^����n�2Mڀ�}|�3�]��")�Z�����7�u����ޕ�=0[��W%1�&n�!������c�cV8Z�����:s����Y��!ro��or)X��(`N�o��0�Y&Of��MZ�qN�C�������m,G�w4�Q���	���!Gs>�3ݓ=~��76�g�s��И�=�U��o���Ã��5ї�L��E���tܧy� &��=��`����F��5^v�����n�(^��1TK�F��o�}��#u����*����ArϩQ!oȩG�.�I�j ؘ�8��u)��Wɂ��D0<��Tڋ<�Z�0w��8��].W,��}�X��um��Ǵ�֑i��Fe^^\
U��?&�
H����4b������-?�")�N��b����R���o�����{�1������z
FW���x�䠉m�J�#߫bI4�ɢ���f�
	�ZgS�5�|Q�~5�%��=M�Eju�W�b.,��]%��:�w��i�!�8��y�f�D�-@��y�l2L�J�~�M�p������Qȕ����� .��8���@�3@zA�-"Хğn�XH�m\u4�Q����*�a]�Ml�ʇ�Z�\<��������6K�Ʀ�+%�P�S`��&?;J���S��d�u����m�J����qO���b��b4B
۟ �� ��ܛ��z������3�����h��0��[#��K�E2���B;�����|wޗRr{|�~�ۑ9�z��3Ƭ����#���~|�v]�o�hb&�IE�{?��D"��aE����`mf߂y+��ލu��S�ʵ�}5kņ}=�Phd�N#��Ff���Ov�ٜ�ͧ��G�Y�?R��f��N;,���(<pܚ���kr�z�Z����?����Y��M ��f�Q���&��� �U9���'� /�qj#�h((K&I�V G��n�vm���S��}���hWME��9ޠa  |a'p��>kR�.��O���t�.�>>���D1��m'���Z�]��?��B�͵�܁���at$M�7'�����2��*��9.xsnF��Pa�'+��7�"T8=��裨/ˎO2��u`��fs#���8SSa���6����.w���	}����f���eg���$\L4��a΅��m����*�z�>���=�n���*J"+���)d��M����U`P�zb�>��v��~����ʺ�}��>}�A�⛑c���{�E����w�M"���/�X�v�_�Y�U���s���Wˋ�
�u:(��&���q�K7�n˒�^���fdVEţg<�! dd@ί=e>;�b``�U��yٱz���'�ms���%7>>$P�-�f���j�gF�>��\�/�C椊���t�YC5 ��7e�6��m<��W�&eߝ���<�'���m�����i�4(�C}"jj>���/>h�Z�:�n='[M��ų�Jp�n�,�*���f�scʋJ��<m�x�re��]�x�X��!���!�5c�=��@x�����_��`��Rsm��S���޵;s��%[�f��� J���aK6�@A���=�,�����6p�%��yX�s:���}0cN����O�7--
�ccszT�@u�q�P�����ٴ�,gF�߳���S��Q�6�G�[p(J5���ȳ�9m˾�d�\��y��ܗ�.[��)M#+��Gр),<]c�����e����U�(t�mJ����}�ŧ���<ER[����p��Os�1�c/����Xm��=CW��Ã�P�5�^l<ؙu~�.|��<#:/����P����8����fQtgk��gv����D���8�������`�Hj1�lqnZN�ZR�1W�Zm���"��|I"!�N]P�E�OY4��~��b�2�!�?E���ֺ�H�2 3X��ރ�����贸
2�����l���d(�8��2��O�q�G�_���m�:B�/GT=�fYH�n��o1����(v�O���Ne2��	v�Ǟ�er�@n��Y�;JH	BI}2�ҢikPwk ��?���S�P�	s��!|�u���wn�;<�KI�
��?��i0��-%X�vM:��������?��<���z<��D��퍎��9:�ܴ�l�;�SfI�D���F���L�v��a|8�K,�:��iWZ�K�o�`V�Kf��h��%�qJ����"����~��:Ӕ�.+kC��\��A�i[*��*\8��BE�0�}&� Z;��֝�UTa������� �_hɔ�08��P��1&.ePT���Y���O�wr�)�OҥY�KR�RRe`^�( �2g)�;�f/��$��O��^L�W!h&H��� 煐(�Z���}4���rS��K��`�	���x�"�DCq/v�~�02_U�G,�Ѫ�YN`���ak!BJ#���)�Rt;������k]�������Y^:>�fX �h���t|��s5ش<沈8e�8��rP����K�O=Iϖ�85.�3�.t�i�	�<��������v���CƖ��/�~�e��gu��̜�#��Y�<��d��Zz킺]����)�3̇$[��3k;_����Y���!J�Q�K5O1��M��q�e3v��U�>��8���-��yGn�uN�D��υ�E`8�
��dj�8�F/x�:nAoJʟ�Ҏ䘒�.�:��Ƈ�c5�jh����X��q��'ץ. c�K�?� ��b�����95%#n��j-	u��V�Ұ�+Q�g��T���|kiA��>�5�ʆ��O�|��s~c몕H����<��4|I��8ʓZ���=s��t�G�	�L	�z�%�$��ᠷ��K6t���;���M"^����s�Θ����]�ͥ�?�����qfY_�u��=�b.!~$O����Bo��!7��hW� �p�l��
l.#1z�"�G���)"�6�s
��"U![���{=5���eUyR�r�?��+U��h��DB�!<���a�|���/x���v%����X�[u�U���N����U#�z�e��'�+!Ƹ���9��XA���ގ�*���}���W��D�5�:q杒#�q�Φ&ӃY����/I��@��[��c+�05�tOM���q�y���i8��	+|@�߮	��	f���)"��kkk�-�/�M�ab�@MpX~x��t�$z�(�G�f�g�棌�(}�Îu9���$L��>f����9E������S�cO<��t��"�(�S��s}ˉȥ#ɺ�`�����U%J�y�#o�Mʃ� �R@���:�R&5�<�z����麬hO]u��$�oK"�����3��c��k�%������1yb�*�G�CWBA���w��z���=o)suu���ZHu'��٫olw��Kٶ�-��o2��E)�����~�v0���;S��ym%4Qc�Œ?r�m��|��ӭ�|!$!�����7�n
�?"�z���,�!���!.$��$���j�.�J�uix8��@�_GLœޡwI�,v�,Z\/vD`��O4"N׃$�Iv��sLw��0��C��?�4�� ������̺be�r����y s����)$M���1%��y6��BPa�;a�}������a�ү�J�^�`��E�#p����z���V�76�̱9T5�\���6��0{��e��H��5E�ddM3�b��F���ri���>��B,�ⰍF��	�������[�^�:c����E9�:�kq�h��r?ry���� �Ϊ�/tl:�5��&�)�`��F�o��9�bq��p������ jT@���ø_q��͘�9�&�\������]�3��Ƞ�����HI��xC,x�x��!P���#�y{'!�~^���Q����<Z��*��;�r�_���t�Qci}V�����˞P�(쀘_s����=K�~��Z)����Q7���RI�����;�+!�9=�	p>߆�BZ�.��ׅ�eo+��n��d���F�U��:�.�11��w�;����~x4?�AT�u.�5��ف>i�aI����ヂ�h��sa[%�t�r�H[��W�]�%	�m����Vb��$�&a(�UTw���e�Urn8��
<}Ϛ�6)!5������%�&o7�%��;�;s|Q]%�C^Ĭ�U�f��;F����zؾ���#�v3�42n� 9�q)đ6��(�0��Wp�;��&l�|������*�<�y^�1 �,�蠗4�������7)��p�9�w��B)5���c��0j_@��(��V��ńu��� 8/�)
����YT���y$)��KM=�mMz��r�B�V�\tDI����<%��i'��@�V�y檜���z��a2�"�.~�<��aS�,n�Z<=����PE��vƶ��dd��o�"�L�蛏i���]=J��>2f��	6���W�;�_<�ij���۬�XsrB�F�m���Q׃����-�������xϋ�c!# �[��O�k��!�^�W�[A���.�":ۃF�� �+�*�~Kr����
���.J��ˀ>\�4�����,�I.D0^ `Tߌ~�DR��%��)pǭ��T}&{�ܶ����؄�&���ڐ"�k�_&8�x%��#�:s�Q$�h�i�k���CV�QC�K����S��m:U훖�jd��<ajƭ����!fneݜF�定�15�'�'�bǔ���)� >����P/������#m��_�;���L�j�I.2ԭ`̟lO��3{<@EMM���r�xF{N���:��՚q���-!�����9��M�~+%�T�W=||�쪝< ��m�_7�̲�e!���а��}S��F��A�B	� ���R�����)��du3��2�yw�֞9ק$��weh�]>Q��[��Lx���{�Fg��An�Up�I�O���h����a�����'ĤHv�}�t��U�f+�sƐz������2�-�vs9�)� �
��O
������*0|ȒH:e9��E!q.c�?��P�\��0�����"7�U`p �f�p�9��t�?L�갟��.C+�u��,���b�cKG��.6�U���9�W�/�6X*���k�4�NL�B%z]=�p�a�Id�[�f��;��J��"�.�$�'��f�:pUsW?�ޑ�N� �|Mn&�ZuO��z,ӵU�	q����:j�aB�G���&�=��^�n�$AM�ğ���i��Ȁ���gql7^�%)�n`�o��H�=�(�wCė���=_yW7�����H9�C���Er#$"����Ԋ����i(�X��6��o�l���Ё=��zf�1���r,L����*���Č�r��L<(U��/S[��>�>q�QI��V%va�}�SKF꛾��$��G���CZ#�(�=\zNX�w�dε7[B5�1�=`��@:�

=�)${/����
���7SU[ܽ�%��W:�g���A��?.�P�����}��o��#]����+�7���)�t�c�*�c��t�)��4[ZE#�2�ƚ�]���4P�Wc6���](;��^���~~ÿY���0-���{�aA�Cqȃ�Sψ��z���.lXDA@@���S�[�D�D�d`hP@J@@��n�����c��?��|����֚5�a�����}]׾��>\�u��Z���Vu�T��u�8������!���+/�������j'ea<���NKuN���S�#7=�̲��V� ��		�C-p<�ʒފ�B��?�aG3hb��������U�=_��}����P�l*!,W��#
$�,o���i@B����L=I�٘�V5_�ϫYU�Ze��*s{�rCq��3���R�gdCKcfw���//VA~�˿i�9�!��>��qc~ dJ�y?��]���U�&������I$�-�@x��[6S��Z6�:cTTԄ���BlJ�(��ar(Z~�*q�rvF�j�a=�4�;X�xxYJ��k��2�V.�,J�$���fDE�$N�.�$��DP;�hŵ3�/~}<�:�ɱ���LgX�}�;&��$��l�+"�\��Q8�.���K�k:[��#>����$�O��R��Mk�������D�A�뫍��!F�H��*��8x�cԂW�x .���y_��GלU����恟f�C'*�g��˽�����=l��C��B����ؼ��l��`�L�& r?�	�S�s$�\k�$�m5S��pui�Io7�˙�5TW��v�&�J�������LE�斥Mf��?^�n���p�]�9��<�V�<8?	+ϧ�ST�U����J��Q��vf�*�Wܒ�P�zȅ��������� :!��i|�p��hy��Z�5��=a1�<_������>k��,�⿄��|o�������N&�z��N��ʯ)�D��L���tq�ϐ^7�^Z���;�u�ퟑFsv�ݯ񪟪\��"����/����hꡖ���'�g���
)|����z������UB ��\<�-�����oa�0�q���U
�m����X�}�d39qo7;�acIr�����X���{����1��]�D�'B�qٗåa�73�C�b`�`���D����~mǡ��������̠vT�YK��t��5S�&Q�K��q��}Z���s'�I��t#=.(���N'�A+�X��S�٩�Sφ%a���F4.>K\�g���˧Uj,'z�1B�H�Ȇ���ug�I|L��G�R��k�{G?�  ꝶD�����ձ�9�ޓ- �]) #��\T:��	�oϮmG��O���.4����8�1����NS�d�:���[��Y�E7�v
�c�ц��,����B��;�/�[W�8�G�;�:Ri��l\%�KRa����w��4x	p4�&q�֭�U����
$)*����6�Ӎ;5�� ��do�94؇9y���q�^��e}�^C�q�f�����E$\T�^
��y�I���̢�gf.*�韇\�vX�a�/!`��J���
�:1� �2+ţ��2�C��znNO�y��s�kf8������H	Z��裫�	��Q̣�=���UU�&~9��	`/�u�h���ck�]���N���-�xA�Q�d�ϒ�	���z{T���Lu�V�pE�ֿrV���ok�!e���Ob#��_�����v�!A�M_w.��	�8�3枙%g��C����m�-�cF�dN(�\?M��7D=�@�e;'��
V���a����`�7�Z��%O��i��{�qv�L�H�1� ǌ>����-�'|�XۣϿZ&L�k��@�ud�ݚ�0 ?�08��W��3�Hw"��6tUM�@V�By�/)D9B��ab��<�*�[�.0� �� �'aM���&�z��K��L�L�VxVh�N*��vŔ?�����m�󥹐o؊��{�'�'������]�O�������w��%}�v����j�l ՝��)� �n�uE��r�ߑ��?nK�Ӣ����Z�a��_�46�@�dr�hS&��:/�D)܆i������O3����CwIy�89�MSe'h�+����*v�������I��@�')j�^���gڴq�`����bҡ�ݩ���K����a|D�(֋d1�7	���a�* �j��DM���l��Av�D	OI~��r��>/���JbA�5�W�ܔ�gA�@J����4�S2�7��YQ�ӝ��LaJ�*g�g��~4?Z$.�U��|�`��{͇%'���U/��>�W�v�?���T�`�ZH�H"Lh�T=����Y��e��f,��VWL��(���9:ύ{��5�n����j�3������M�W��(�	�ff�te*�z�e������Wh�C7�CPz�{�D�+���׾1A��`n�"��[��<Jsח���xw�/�X�r�IU��4�i���N�8#'\W�J^9Y��1FK�Z��<�7�P\e.>,��g�a��?��M��I%���cv�|^����,����%���T��#a'����ka�{��~���s���Rf�K�����J?��q��#��
¥e������!��x��eg����8��LW�.W�(	�FU��5��3�K���*`Y�g���޵�J	湸��>��ez@X=1��>n�����Zŀ�0�ڃh���?�e����, �^���u�Չ/F�(���i�q �MO*Ĵ���2�r�j���j�@���
�}��k��� &�ﲷyr�KI{T�M�Rg>+��y�C�)'�Ѽ;Odǉ��LN���m�P"�D��a���X�ϲ#�tZ�	E�c6�%��w��?Y�R?�k�����G�����`uv�e+���8T�-7eV���,�K�R���c��$#��)Y�L:��m��NK�#�f���k�;G,Օ��*�o'���29HԶ��^�@>��\�)����N���#yW240R�'k�B����ym��ƟqJ�+��?����-�_�,6��]��>�����3�Z;:[b�~������aWr�t3�=��r&����ԋo�Rj���ݥ}���4��¾/ofo�D��G�|n�l
�a[Ź��ݬv�7��x.f7�vȢO����LU��K�	STL�dmfA�C��+rȖO<�*����l-:���c�f�%�QPb�0�}���fZ��F%����}3h��V��K0�t;%�-L;�E��� JM�M�4࿧4@��h8���Iq�?��ɑd�������!��;���3��o��r�Ӱ�!�cMr�.b^R0�;m��q`���~Ba�,[�g��JKѸ'�̺8�
�7�����m��p�w)��?E�ΌÍn�p�>-�����|��[֧�@�W�xJY��q���z����F�WX�@�Ym�e582�J��s�7��{�y���*q� ~vQv#�li����b�7�K
,�abwW^(�D>L�������������u� ճ���Ez;�F[�K�1F+�4b2��iiAU,ݹϧs�.���F)�1�
�x[a Uя_H0��+p�@�/������N�[/x�����
Z�ֻH�@�8�o� /Ltw�C���ծH�M)�����'�:�	�$��d�/�3 �H7� 4D�vTQs�M9��Hs���2�z_i�-�gFb!���d��O��2��P����=}�z�oFh�b�]2�ﾪf.	93�>�����b(y�ғ�*,�RF}sв�>������-�{Rϻ�-�#ذf(�}d�2&ל�s3��_�D�����K�%���y�A2<z,�o�1�D����Y�/e�eA2<db�=�gu����|�οظq������T��/.�E4�֔1v�kiV��eD�I_�� ���A�M��p���"�'��-��*����Y�d���N�� K�3���ܾI�i��v鰏%>�Z_���?19<���!,��㲜@���y�s���
M#F��7��_��2�+�NT�͉��8*�5s�ι�}+f�0�r�R>���-��������D]*O1�F��f�Fj	�I{_��A�C5���\��ɭ˴߮�w~�֕J>Oؤ�>1��%��<e�4��O���?+��tV��c����� Տ[}������YC�e���}�T�W�n,��w�AmR�j���<����Iҗ�A��=D�G:�a�a�c����Nʧ�=���l�a$�!�����Y�L%�8� �O}�Â>�+:�F3L^収?;��ev��H���_=��Ind�O�mr^�v=s1�뫰��p-��M�Xő%�F�t��y׃cY��aY��O�}��� �E6b�G����A�5�d� A����M�_�fw�2R�9�_Kk�{�:���5Y�������U��R��!y%^
@��36���6y42��̃v�(JU�l�[0���B�5���y�R�G������)տ�,�?�GXZ��4�G��|�촌��������!3#���p����A����],y܏ |���Z�G)Dg+��͔r�1��gvw��ر�G�unu�D�B��������hƊU���`J�J2<�؛U�9���]*�Q]�sw1Ox�|�����tSm��Ʊ�,���
�3��a�Ȗ�K�ڣc���U�7�!�?B;��*���tvX��ې����W>��F�nN�ŠN��������ytx =�IM̀��"p����-�?h`��mJI8�1@�<9&����)�~�ظLǌY�$���3}�#Xq�Q����LU����,%�x��a�`ύ����:�s�z֬�k~E��p:��d*)�`�AM�i�xBm���
L�a*����~6��l� Sˇ���� 1{�M�Zj5���F#�+���*nulFw�ƛ�����H���� ��r��L󣏖I�kqm�w�7?���^�[��̡e
o����;LPLi�oG�@�ڛ���&���N����gR�vN�Z{.����� `�g����?�c�?���Y�Σ�jM�x��y���JD�fZQB�y?�9��B��F��S{��߮�����j0�J����dn�$o�W:�kw��"�B��Rq�&n�Ҙ�{��&JT�� ��|�CS��)*��H���._:h� *��5f���"@�\h�"��M����8|����˷b9r�v��+��"�:%��^�r����	�\�(�������,�t&���z �j7�r��$ڤ�b|L|�~�������LB!aN	�z]JPm�s�h��x�]m�S
��cG�W�ҳ��?�+��:�����&���8����R�4?ِ�uNqJ��~z�i�P[#O����n������v�ܦ@����.��Ô�4Y�����d��U�t�d���[�:*�Ѹ��v����Z��=մKDIj��+ZHi�˅^��
e��-7?8;;����U�Zw����cK�Er/�#��E���;<MF������k�<
4��ܕ�sC<E-����RL����K����F笧�4:^�zza>)��̏#�oɴ{�X̐ikj�b�����io}���ύ��Q��b����9�0����P���+7���t|+[rD9�64/�C׉oOlw�}_T�Rg,-[��p�9�<��g�d�+>�Ķ0�#��N�A��40��v�ދ���Y��F��s�S7�d���nߕe�Yƽ���}�d�)
ox[�6�o��c_7�3P`!�+����k�B�m|#�I�|����W��e���|� Z�S���Px�	�f�a�0����'��;��joD}�4LE�	i��Tf�p����hX�!������}�<��;�[2<�=q�I���e��x��Q���&�Y�U���Ȟ\ncd4����*�����^t��|����:`B��]Je���Z�$�*��/����ՆӁ�g�K��&�]]<���ˊ�--#\o;�7���&ja���u,�f'_��#�Ϯh����.x��������������L��,��tN���b}�iWN-`�lzB�n��~����E�j��b�P?�Ι��.��OW$y��!�^o��{ܵb+WY��K���V�5�� ��k�)Ka��΀���� j䕳'�C�zB�]�K[W�-�H���A��)�tXa�ȷ��N-d�%�J�ؑ���O�b�6'�@��D�U��	j*���v9�<�5.�	��K̐o�.����-�����Y3F;�CaYJ��o��e���;�&���7���>N�)�@�[�ע�ʜ�;�J�t�[��
�:d��>��{�I��>Ȯ�.[
Knۛ9����X�� �����ج���v�t�-T-_YĽ��Ut��~�fw<@���;
ø��
׿3�.7~�}~��u�7+�A��W�K�f���E��'evb�z���DF?Ye�_=��#a.��[4�a�;�3W;d9vO���k5&�NRNC�o@7�3�;��asj��������ڛ��~�����V*���I>�u��g��)��Ll�;�h�:��u��oY��z&RL���;�ø�ӆ�'5��4�NkL���h�0���gY{Rc�C=${�DK��p#�!	�޷8nb륄ֶ�_�FIZ���i��P��e�KG�.��j9B3��"�ګ�o�攴`n�2�P7�=Q�����Y��Ҡ2�n~��dwس�6�bY��3U�FX5>T��ǟ\H�m"��0_��CV�A�=Ƕv8�a틍'W�d�/�i��7�_�(I<r�6W2l�I{�yB�O��\�Ҫ<t�.]$m�9��~�J���Gz�C�H���F{IO��=��2P6^�ɤ�9�A0А�*�!-M
����޵��?� !�YI�{��f�U���p�ulJ�Tȶ�]N����x=G\�1[/.xK�ˢ�>y���NS0�%�)��O��c��r|d�������X�!�5�(���s��Kj����}�h=͠��[��5Z�+���w@D6���l���qHj,W�M�V���u�x&�/�x����~-0S���Kz-��T������N�����t5���&�j��W����2O^jp�w~�_�8�m"�t�Z��C����1r��^+�Z�VtaӸ�lԉ�Z۵�$��D��S����7HED���Im��<N��'M#��\�#]�U�|����	�:��e)�)Pp�M*A+�$G$�"��	}�~ja���2�d��
?������m�@1/O!�3�bҩG��a���b���R`�ֲQ1���%tDs�����Ki@�u�d�k�n�xQρ��`���a���0�Y�������a���t�}�x�1���ʌ�
��*�~��?�W/Ϣ�An>웮��g�D!.!H9aG��_6�`��
��,7<���z��i&�{�����zZ� ����ŉ�����Ҽ"D�.]�zc#yG<�,a��z�����x@�i9/�('��A���2h���a���Jɕ ��,��"�{��A��l���s�[tA�+BjǃY�pNԣ�0W�G�f�$�{����ߌ� �:,�4cC{�K&�lz.���%<��n�C+f��k)���:}Z�^8�:F�����CY�J�q���<S��w�����I����4E� �8#5&�Z����E�t$"E���P;=�q�<�� o���ă��3�
o����eAYg%?<O
'J�[J�3�n����
M�4˒����3U���O�,�iٙ���v�?]�B��}�c���Y�?�p�ԗ��UJ��6�`,�=kˊ��C�6j��e,�u���y[���ȣ�[֪d�w�cs_^'��eM����ia%��՚qpc�:͘��p����`W:�t#i�����@
j��h�u����C�F��(�{�֙�6��ɸz�|���B����a.I�j6J�_��|I~��U7�`��E���*p+�ퟠ��5���Y�RLzj���7�@��K=���ٳ0�qױ�4��X�
�B�������?0@+��J&�F�W��܂1�X�� "8�\.�Ʌ��>^R7af�̨�
����]��~����T��ـ��K�	���Uy���}��]�x�u&PS��FDVivZ �uJ�?���E_�� (�w�'4�03����|��,F}������L�rk��?�Z/���g|�S��2,���Y��=i��Xe�=��G����̯��-b�����"�g�/b�f�Ee��B6�g��#.K�(���B�lG�b��7�UV�,B��ܥ�Q���ݔt���=��7��������h��Ւ���ߋ�7@ �Q�}2� q3~��~���KB]U�q�?T:z��1�ao%�I"��TF���Ό{���	����s"��b�3%I������!F@mpbȾ3��Ikwt$I��W�������xz��}M���R7��S���B��l��@B�/�l������X�s$����4o��0����������0¸���ͨ���ER+�{j�����qL�1xѠ�|(c.�{�=���1~�G0VV��ɩ���FBT8�jޱ���>rt#�X�����c�=�Ҫ��,m�ԛ��OFA ys{-J�Z���r
(�Ek��~�l=I�Zi)��W|�H�b JbKN@ڶ���XsC�*܋ޫ�1�_��[���O�
�O�gLm�A�<UKc��h��l^���
�g]Ӕ����?�$�^s	U|NG��Z��>$�5�I�����5b4��������\b�d���$Lq0������.!Lk0|�lD�ѐp!Oc��K�~_�{D=M�L�����R) �����LR+�������<�{��0��kP�V��] &:^��umGC�3r������Ȟ��w��zb�E�4]��~ �?��a$���bG���+��.�yx/��WwE� �V�j�NW�=��9ߍ�W��o���۹ā:Yy�� };����jv����Yf��h���D�����n�bAC����٘�0B���F+��QD@�d�4��:�ykX� ����S�l�M]������m���}�H!e��̑�"Rd��c��#�vc��cCq��5�Qc!B���J��F�)��<���-�����~x��u�=���J�MM� P�{���[�G1��3$y�� �.����>�E��(_Y����v9���N \-� �$1�����7�L
k5uܺ�/���$"�Ne��F�=,7���3��I�d����R���#�߲n����p�g����l����Ѫ�C�Zl�(����ʞ)����~�;����E߫��|�n��t��Q�+���.kl���D�Թ��Rz����1���upYu	��X;@��إ9���nd�=�<�8&g���(���'�%�a�ҪbK���H@�����t���p��%左�za뾓��F�>X#,U>:1��,���&O:��C�*�Թ�i���������3g
[��p��.��8�k�������X^}dfl���R���<q,v�\-��@�(������������>�c�V�@�M�k��A ��#߷w㛾��Q4���+	uB�W��Dw����y��O������oc̥�p� e1�cU���2Kp®;bћ6��k�h��֎��Q&��s�D 8*���DMӖ�"�QC�ߠ6�Q7��o�1�� �F������Kq�G��GmrT���d�L>jY�GtTj|c��6�.�EP���^��0�b�U%���_�ƚ�iHY���x���� �� �4u��}�ʳ�\�Qp�s��'���#ٜ�>�;i���|��y�>��2������,��e.�ï(&��"�i��(����5v��u�����]��� �zc�u�o�nh��2�F55�ZҎ*���N$ꬷ����SҜ/|m1����I���~0W��9%/���������I���4�`�h���g/Ŕ��=zKP�f�Y��S�'&�6�:ab��Wll����N�2�ND�.4(I�ʳ�v-�NP��-�?���XS5���ǃ�6(��M�|�Q'�6��$�J�P�6�+cxk��Rh���w&���Bΰ�������/�~�#�'����&A����l�0M�CD����7^�,��1;����(%]J�dN��
	K���w��)n���%z�?��ŕ]����oxh�3�i3,���]�Ҵ��K%6B��<����82{d(b��j�qP�T�AF��N��VQN���'VJ��?=*D�$yyG�_�.�8v�2cQq �'n6��g�I�N0�}�q,�?Ʒw��1A��k�F�ly�@��ZG����jޢ��ڈ�?G��T��ΑeJ�O��=��M�L��?~�H��?@-��5�砕�L&�;�=�"F�dҋ�w�B&�%xG3ކ�NZ:�_9�Gif����;]$a
E���>��Y�(�*"���p?�Hy�԰�p߉dv�0b$@�_�ŕ��[���U$φ@6d�G$���ўN(��Ƥ7_i��
�;�t��(�[K�@c� �v+�"T�'k���C���E��	��o�ҥ�n�n���0����Q�]�k��~��2N*��y�-��Z�8�8�Ɲ��?�	I�im�����}����ߋ�tW���H���p1f�  �͋5���}�֍��[v�kKZ�7��&����ν+]���Ͼ��`2qJ��0��Q%w��ѐ��R���0b`����ͮMd'3��}���w­�CQpŀQ{|�k�:Z��;<����	�_}�~���Ƒ�4!���_f>3[(4�5��cb�3k�s�K_k�M�M\����'��F�2��%�,(��̛�TS؊6��^2��ꐅR�J�hW0!$�['��-+��E��{@J�>�����p�BY����|�9��a~tB��AR����입\�5�'Ի`�P���]\����8s$��ތ�����\�hkb�/��ͺ�3xRS�[A��\�	��gfV��?S
?��������O��(�9���{̜ɇ.q{0����Qw)s�:�g�	7F\4u��+���>ľ>f��)..j{Fn�"�Eu�c �����RB�)�D�v�R^A�r�D(�8����/�l8��<HRƭӋ�Q�N�����k}�����P�o+4H��r5��V09�}R�m�Ra����Bv�6� �pe��gGp��{��y{6|6f{;KI�R��>�.��Iw����Dg�T���a��(�i��e�Q�挲��/�3�7�do��.1�͎-P��wY���	��s.v�1/��	�׎����W�a�ũ{�{���{^�ںۯMzx��V|��f�-ݳ+D�?u���RӮF���?^��֯���z1��o�L�Wq�M��́��ף��9�d���\싶?I7J�ҭ�4O��6
���+��S�$�2���������3埭q���ߊI�ޞ�
ܢ|n�oT�Bm�6®]�����hZ^rw���#۴!�ȫ-�������)��+�p��:q;�&;��j�(�4�;�ţ��@���f�DH�����x�>�R�r2�$�~"�P����C0B�J�4�&vT�
>4B������:���G�y�FeQ��W2���(���%rqS�w6�;6��]Rէ�����Mh?L�j��6W�����P�Th����O|�C�2Fė�f��V���	�QV�����F�G�[�Jy��y[3��-Ȼ���?��N��r�e}a�Wsԍ���#hb3�� ��'����$o6/~6�/T�毹,lm�f�T�۽m��UG�����arI�9�I�ӑw��.��qф�ඓ@��o(tM䈨� �4KL�v	�7��	S�{���ܚ��y�A�OG�b�n�[��Mه�����0@����W��9��5��[EU'gn���,�o�'�eU��*��|oj�gr��������~MZ�YD8@���W�ǳ��Y
l��� `�u�"W0*2�6��2.��_Ǟ��yO~��������8�nV����n�i�L_��L:��␢��פ[1�����lu���wSwzx�}c��69P6��J%�L�8a��	z7 d��5�~'y�N%O6�'�p[P�:�*��B8�vL�6Yn-�I7�T�u�:Ex7[TL��\��Bo��
�t�JZ_8���j2�+>�9��$�J��Et�a2�$��@s���-���2�	v,��}PO���.5�̅�X�XR/��/g��VzYP�ye�-��}yl�.@��B�\[_��G�R�L5�{�<��[��i�<=���y�m�7�4�[�6�[s4 u�Ng���5�[�wDhmU5t�*�v���L��{�ee��]�ȷ3ȕ=g�ZD��_	���jx��p�d����"[?O�ܘ���O+�9���G���U�]������my�K��9������D�QFm��NxyC��,�rk����u_�Yw�q���n�U%@��7}l��_�Q���K�ں:��V�،n�u�ȡ�h���(˽{�d�4>��w�(��Y�ֳ7�.��Y���|.HUl��a��V�խdA�P�Sm��	����L�Q����
W�y�6|B��v�i+w���;v PD�������o�ڦ�����JH��P9��ͣ��@�ml2�w-EJ�'>�p��i�T��K���1/�9�!� R�� Vz��¨^��0d{{Ga��°�r&á@��w�x���}P@��P�����sRֈ�[k����U�ơ��>���2n����9ݪ���Y��P��|�{�����x �S�ɼ��&�-Y|#(���R��y�E�gM�j�)-��B�a�P�n��n��~,���u�!�*4WlwV�q�/���Q;iE�u@&ؽ�^��[!�q;W�+F����F�a��	����aB���$�Ӏ�㠅�Q�_����j��7@ 3 �nR9�������A��]���#�o�k��{����h?f���
���}���Ө�H�	��6��tZ^zZ�8�ۙ����Oe1T����c3������O
/�e��׵o9l�"i���n�י�gmX���"KȩqeS0G	-�ڔ��e"eou-P��%mӓ�Xk��=�0���f1��cVe+��3�y�n=�����?khMq��V��s�86�/}���T[����K��6��d��wa�wađA��n_�����#���Q_@:�7,`4��x����Y:.x5KO޺@���Q95|��;� <����ݾ�ys|b5��zD|`f�3+��	�(jN`^*>����!­>���8�6�"d�y1��i]���>;�ύ{�9GJ��*P����n��1+$U�@@�8��0����V�M�x����ހ�H�#:��c/DZ}Wq�y��� x/$��������U�����5L;���SA;��俅��$\;˿��*�b��$z��~0�F��f��B|�y�}cR&%��:� ����$���R�{�%���6���m��9�����q않�����KR����TC�>ݛ��1�մ��ʠ[e��.�z��
�L�ƛ���Mĸ��<���tkT�g��髉)�l���Z!�0�r4�u�L�
��Nn�3�Ye3�?~��.��vÌi��kz�
�p�YvL���9�U*lI�-2`T|�P�z,������۠��g�Ac���>����x�m�{�~��L-���<�c�K6��h�!0B���L"l٪��*�Ei�.nR��h�������������I�x�К���:���q/Gq-��/)�q��Ї�+�B�.�[H��#�1лP
�Me��QV)�\��d�
�a��8��[9y�{:k��͘R��<g��yb���K�^U�H����Z����y<��.�P��{f�o^��s�~|���u/�~�F3n�\�=���N!$��\u�Y���� �T��+�<G N[̃��C;q{����y��l���Ak�4����&ų��o���#䠎Y!&��.�Wޝ�
����isM-Ƃ�*��nN��u�3��s�V�G/��6�"vR��1�A]z|��g�m�oȼ�9��:nyC��EL���@�U��iR]\�8ؼ�~ ���b�Ɨd�Sy��_=�;37��v�'=��=k�U%E��)�De�~�,DLRh3�
��f��A��=]C�*��a�Q���rz�p�{�Z�p
Tz��[z��!�mmE"�r�&���ɸ#�l����p�$������ɬ���,���G+���?��76����1F;Q��9Lނ�xl7��{���xzn�8f��VFf�����X���U:p�Q�A��Ȍ���4�_#�y!� x�Dܮv�Ǩ�whR�
g#�V!�<�Em����a���m�I�Y����a.����v��aZ� ��)�I���q�%-h;e��Fj?)��5���+.��M�vu_����Ҡ������̞���X�a�AiX��ݝ�T} UV�7�a�Za��&���z �߹C��vi�԰����k�9��'���.mq}íct�)���VG�9x��Q*q3�l�]��jL J��G;GZ�	��f�����e��O�,�y���xO�+O�hx�ژ.;�[q�*����#rF��2%jf^a[D�w׺4Nw�W����\��Eeaa����y�U�{)��}��z���貳y���xs,�^�µ�����u&�(a��"D�W��-/��)��	$DZ�"[�|��i�����la�R&���o��
��VRX!�ҡ,��~��JM�N� d�j�<ލ���2v`��6-gp���L�5�y_ի����kn�!��V�]�n#w�G�k�Ľ��4�X"��O��(�]b�2�#;=��ǎ�b�a޸��!R�`�RM9��F�R�z+�»'����>3�}�4s}��+��ă���Ԭnnj�����&2`f?��dՂ;��v��sg�V�����6�}������%">G�\u��@N�V���]ڷ�ۮ���&�ʿxT��������.���@��gE��~�Nk6�ۉ���xUڹ!�~�w�(#*=�(�7մIEM�yk�~�V�B�)���ֈ)<��/ﺇ��1T?�@7[�����|x��@K��;�'i�&�a�nM�
_k�SO��4抩)8*k����g�nyp�3�4��.��4��9����BT�ۼ7zD
���D!`,���3Em ��+\�q��w%�d�&�m���*�/� ��PO�� �`���Ѓk�!L��=0�8zGV,�G�n�a���a'���D���5��*�zC:�^-9S�l_�ȿU1g+-�-/��܄4�Ȧ��Q)�&�7��
m7���������L4�0-�P���ޭ����� <6��a�d�C��v�n{�C�P�
�=4��N3{�m�4�H?��	�{tz����;�Ba]�(��W|� �4*p�� u^��]�Z�׎�/��¹�����7Ą���XŰݠh����_�N�� �`���Q�.��>�x1eT={SA��������\�U:@;�k2�	��,셧�	3����l��k�'��y�<��YNt����{� ���jNjɿ{E���=�얫�ʲ�9�n������Z�e��k"#��tE	�\ݎ�L�� ?�3����dk.��2�ħ�&�R�u�u�й�M��(��ƿk�E���<_�Ќ,��۷+e;��N6f�����S�yl[�99z<?<~һ��9��kN�0�rXr��f&�26���hŎ\;o�7F����!�A�p�O�I֧��=���6H�T̆���� ���:٬pכp~���o�RD�6�9�K���#$b���j}8q��Q��E�7��f{IE���*m�t��ǘ�V.��d��y���E�J����
����	}��O�&[/_v:��F�����n���)�&B�E�s��7��Y���:�`;�K/@�E3f�j8�8,��"�[\3�F�@=ke��@8����8v��d���"ȜOJb�Q���ٽ�N>]rA%:_t�����fx���$``�}a&B秘�	�A�����L�"�J)nYE���ws��tr9���o�H��Z����m��*b��ښz ��V���������L���Jr<;�ħvZ��S3�h��cox2���f����P��8[���HpD�9Ӿ�(�{�ҵ�=�&��Ēۄ���gq�s�Ө�|I�K�&G��$�����.Ѫ��ݟC� �A/Uu��fp}J���g��[���"c�%�baq[��w+���#��I���x����7��ª6�s���ޕ�Dě�c�J�*��n*�d8��>�p'�L�y��������F��Q�M	���
od�BNLֵp?j��Dy�����hjWt�̀�&���m�HLs����#MB� Q"��BL� 9"e\v���ջ�Ν�#�7M����=�V���qS¤��Й׶�����.۾��s��j�+�o��Ć����6vN�G��l�?���u|.k��PRQ��M@��Ae}��������E{q��K
����ƣ��&&�JJF?�z_Ś��
��߄չH������Ø��szF|^@�l�j��u�����yV�-ٿ"zs�Υw�C���JM�O��u�<da�r�}mj^P*z,���$��GQbM��r��76
��+�k���Cע9�拋G���r���&�>�b-t9��!�f' '�G����7z��:�V���jE�/!����=�5]�bc�3��l�VkeUpM��O-���+,[��$R2����R��v���*�[���ۯ
X���
�.bߍ�z�￧s�+"2�~�(❷�W����z��o��T�d�P���V8���\�V�N�$�n��8-J>Rn�i֮U_��)~7���cT����C�3
�0���X@ c�s���䆟b� �o;���h�s~�J�>�[x�e�La�i�c L]E�}�����{G5�u�Q��Y�-�H�#]:�j�)UzWB�	���M:��� ��J��[h�J�p���~�;�;�=㌓12�h��,Ϝ�y�z����MZ����,0�񠜖G.`ʡ鹽������}�g��g��"�LQ�
5-[��aF�Z��vp��q�uxz����;�B�2��5k٥͟2�o'�!����8D~n+�P'݀��5���c����_���O�N<6�35�hv21z鉔���ؒ��mN~���f�Q���!�4���vת7���c�O�!�ͽK
���ό���6�.k�(&IHxm����M���-(��S6&�����ՠ�v� ����,4I��
��0���qЭr[0���s�#F���q��ژE��L��Q4Pa�����b��g�&�>��[����,!�����'*��n@�K"�#�{�\�#E�Q�=l�B\���Q�U�ςK������C�lj*�L�.yk�����M�	����"ǻ�EK���A"7E3�bKNInmP��=dٓ�O�1����Ј$��Y�Q�l�	���[)$M�/����Z��g��vlzrV=͙J�i��x�,>��Q�F��E�|cRq�M�D����}d������X��o��Z����2��lR�b�gZ��b:�B�yD�������"�L\�b3�m���<dǺ|g�0�$�E5��2�&�S�?WT�=n�8BȖ���/	���XW�M�5�LQ�j������K��p�^�oI(a>��G$���D�7��Ǒ�V��4�4�	�H5f녌��:%�����	̹�Ug�6�A��y�h���򥫶�\F���8��ښ�Ι�/ݣeӆ��@ꂶ&�,�4��v�=�c��s�؋�Tvםb	�}�S�2IB¡�o�O��2*mQ���3ffajT�"�{��)�	�8��̕�꧉z'/����	�b���t���t���L]|*��d����-e��˖� Ex�&ս���nؿ#���x��BC޾O�k	��ur�����l�x3Y� �Q+lbiawD���`��(�T_�M�s!U���͘/4���Y��fh�Q�J�&X����~�0/�?X�����O?������y��	� 8���ʽJ���1�ܬ9��G(�XZ���I_P�7%�*jjr��l-?�7�����W�O�Lѭ'��k��YaL;	�����ڮd���O����h�0����Asa9������?�2�����w��":Q�b�Fb���G��tT]�/xl�!�����s��O*�Fx�����~�c͖���)����Cc���k/щl�H$~��ô����ҋR�Ts|>�N�_@��ii:�=�J��/Gس;�o,��z�+I�SL ����c3�.�t�]�k�>KE�
!BCo�Ѡ����	*����%I9�?Fi+]uǕ�.
���qf�������ڸK�� 5B���u�Ĥ�	ӇqO�.��퇊<W�'�|�^!��g��75mthB�:�����਼����#��B�˵k�W�ʖ��F�Ћ�R�F��[N�����,�
��Yh$,�s�^�P���3��:7�zW?�싡r.�i;������:�|�;�h��FPk���A����|�;�����2;�u�Ȱ����C����ܳ"t�ֺ����C�:)�m(ܼ6��9��Ĵǧz���<>fl������:$U�I��Vb��4g���%���p3S4_;�8PN��X���g_&�6S��lc��X���C{{�{�}	�E�x���Y-)�4|�'��0S`�
��K���xH�<�%Or��s8�� 7�[��tX��bT`1"������-�l��*Vܹ�DZ�=z<Gu��(s�Z�4{�甯iG#��|#a��8ޣțGE8���9��L>�g h�����?EG]���7�_f;�L���u��pN��oG�������Z�o��B�EW�fT�nj�K+��vJ�:��/#3E����)	���	�&��o�����<WL�7��r�t���M�=�(m�W���������kU�`�ѕ{m�Y?�[y�Ŝ�Z�[}��F������V#��ֺƈ�z��gOY�`6����BPnO�L��3�^���Dp)V�93vY�}�>.����@@���jȭ�-�hV�A�2,�Ň��=���O�����=d��7�pD49�5��~�S����������斳]#�b��\KNV�u��HC,g����T��6U#]�%*�ʹ��^��!�D'*qg�NТ$�D����z/�!�c���[�OzD�
���^-ұ^��w��,�v(�@;|�yY`kՉ�������6fX�v��$�λuI�.;=mނ�9T�ѣЖb�D��=�[Ȃ�6g����q>Ŋ�(ӫ
�hf�ց��DQ�Ѱ�{{o<��9���=���f~*n�D�C}������h���9NI�����$�##qUȄ��;�)q���h�A`|�/]���V�� �+"�Z�1»g<�7+0�u*1�7�����<�ˍ��ա{�=Eb�[�����Ң���.O���l� �*L���:������V���"3�+�~t�k4�#23s���� ��_��������耒� ��c��`W�,�H8��2�x��!st4�+So�+~�<��#�py](�����(K�5��NK&)�.��9l�Q9�8��O�73#�T�^���*2�*+w�Y�Jt^<+�xF���kdx\�wn��c�u��{C7���cV����)�!I���XE�|Q
<[����EKs*���������Th��U���q��NB"s��2��P�퐽�Z7Dn��	�v?���*�~���X�^��R�7�"��A:P2`�=w�?cwy)�A�PMucfT������)'�gN��\�ϝx���m��ls�u�H�u^�`L�V3�'���r�)�CF�?x>�Jl�"�z���Ō>�4��ZWc܏4,%f�������~���ѷǗ֯!�L7`�z�#�u���o�!�$�?ʴ@��(_��y�\+����L�#�V�oGC�/ߝ�$%P�����ld:m�ҊeF�:[W��J�I[cC�;!߿�d���7��z�%#4�u��s]n�zS�)%�����!��d��r��Us�@&_�EO��~l J�a�pd.��:F���y������&�.��	(���i#��Ԝ�$n�����=����[�����P�1�L�PX,u�O�V2�H�%��.+o�1����\�B�Zw��Jt����L��B��F���ƚQ�aX*�d���_k�M\�M>Tڴ�"4��:�mP�c�����_.]�\eQ������A�ts�&�o�d;jLga9	�\��>�b9��Lֶ4�Jg'O�W�<P���8(S�K��d�H;vʡJ1�� �yؤ=�r�˕$�Ŀ����0�G��>VW5*��ۗIB�r㸱�K97�?�&:����^ Ħ�h��o����7�E۳Lk���͎��#� ��T�W�[y�y}�j[|$�4���;m[�����N�)��b��"��*_�6W�qf��&�N�<�^������; ��XND�@��tK�����Eq���?Ǥj�Ǐdx���N��a����kU�.f&���:�Y��.�6~@���PF7�/'M��G?iX�s��%h���*�n#�(19��wX�B,�0����J쭂��AM�[�i��Bȝ�99�0���)�CGQ�h����G�Sj�T̼Q�0ÉW��w]���Ff��F^E���~�R�V+σ�G���葃ھ��|@DW����Ն�k���/銶���,�´��Ŝ��/Id?4R'��pn��o�]����s[&&c����&t�����T��sv,)�:�:ĳ�q�'�[�'���4U�����0��g-����sҾdf�[AG���g��]�̍{�ڦ����c9-�M��\]jrM�3�z`=p����_z�8��B�ɳ�h�+�\���G@��+X8ZM&�����:@��<��(�m�x�_�������$vG�:X��$�y(�4���2%����]�j6QȺ�c����9�3'%��t���@s���jF�ӵ���o�iB}�F�����u�U����j�md08#	#�Ԍ����t��%gE�D�rx�9i%�(��[՟*=���V��n�}�\��5GB�:����J0SG����gp���!ƀ�'��
�����A��yc��ŋ���DI��$v���4�c:�Sԫ�}}�W���a��0�������.tO��V���pn!�w�κ�FQ��"6��$�KY!�ysl����_���r1^�[K4M�0�6�-������x����c/�Y�ùɬ�6����e2R'������9mJ�ݷ�QTMN�=����}�ﴷ�Ѩymڂ�_�=[�Xx������w��y�"%?��b�T�P9�I�q@J�V�uGJ���X���^����yOz1I��>.,�=l��:F��K/�s���7�m�#"�����1��ߗb_ M<�L_V�G��*�ε�̡��}���ɐ���W�u���n`�F�/?�,�1�3����13���511�����ǐ8^�J�([O���ٷ埵�5��t8fe~%�j���!i�S~Oy��]g��W�V�(�d*��S��$�(w����m�x�5�P�a�O
��J��k���R�8XnX��6$hpD�m%+P��T�u������2c�4L�zVV�c���8\}�����w!�UO�кy�RjVê#��4��b� �2L�C'��tZoU������śƻ���Ֆ9����E��ME�w�d��S��K��#e,c��ɷ|W�Я�=�W�?,j.n�o!�@.��%.�{����!���͐�x5�:V�W��[%nCŅ��:�q>sQ���Z�8�y|]�x]e��=�m:�)I��:�n������RTj�v��m��F�^�����"�9���h�/�M�3�jR���4a�lw��8kt�5�86C��#���[��V|��?�2�ݜ��P���)�mЋ��S��Nq�|��r�GnYn�2�W��i��U����$F��#�y�i�OOO�d���[k�����k��fq�nf3t��S��H�B0#�|��	�0�~�F�8��N�>y&�̓�*���r$k��F)���
H����y����u�o�\�Մb�Q�l����ߘ��������V������� $Fg�<\�-m�| �Q`KnۙG�ai�)�?�u�z�,eec��zc�"��D.zUs@�5��h�5���c�mq]%��P��|��d�#�:3N�9�\��g�J#G���u���@G�x�B4�as�bV�����
ɬ�Q/��Ԣ_/�[�%���ɖ����2�zJ �j����\u���\��Ź��i�+q%�:�%�Y���?�:̜q%o|o�ƺik~&3�K�,��|��㬗niW�躱�g�����X�T��w��T3���� (�:��j���������p�歕%�)���x����EU�؀oߍ�r+���}~��|���58�&��*�#�r��ߐ\(
96�7Z�9Z��3s�� �`5��[��+��k���n�ےf�G�Ȟ��ėS�
���DUFE�NɌk��^�^x���?�;�H �U"pխ|������,�J���7J�5˰����;0ڟ�;=�"I�W�# �;�ż�bۂc�HCVO����y�z�����y�5N�H�!j2��o�^��(�-3�M$��ғ�����b��+�v�h��n����u��֣���N�|�2m�t�g�Q`e���]�b����H�g�Z9Y����!Y��XֹM�o�iЭ�TP펯�_l`��
��l�l+B��q~���ىOR�mH3�RZW�WU�W���x�r+���+�#�Ϭ�nq�}���P�rUx���}�Z��Y��Ӿ���*��;�@�1�繢x&]��uO7��7���fu����"�����l��Ap��9ށP��X��+|��n��40;a�ף!�=~������/Q_1_���B���5ҋl����}��6׵�oJ��)w��l���g��Ew�(���Q�D~������T�y��5,����C�cI�;E��]C|����sf�'���Y��3��0�y�(1��HN��s/���.٨���S�w�P�Gn�\��yge�;�!Z�=C�$q������X��o�M�����GXֆ����GY�󜄃P�Bq�*N�D�sؐ�_Z�~��GQt�Ⱥ��o	r�0�:�
�qr{;G�j*o�Fd��m��_��]v6�0c(�{�.�bضV�b�ڬ6�9��~3��m��.p`��������W��9�y=ƚ�E�_O��6��+h�^�`�8�c��%���k���uc9X1��a���5K�΁r��`�����hϗ�6�_=!�1y�G֊Y��a� PW߅)g��~�_����e]��7q>��=Օ%���v�`kQ�Z�1-���-�}VQ�kn}Ͳ�)/�e-T�̈�U��p� Wd\l)���	�Q=�j�;�p��1݌�>�Ǖ�~��v��w�{�����y��q�9�6u�21���+\˼W�EW���{Q?&�q�ZY� C���zp����Ĥ؈d�O�yψF�u�g�U�=�a-A���#�ޢw���q4�j]�"��Z�����zm!^�U�V�e�н���X�7LI5v!g�yl�eԙ��ۂ�2��75�rl{�q�Y^�l�;��A����x*���*4����.�}�^��,::�nw�ӰԃU淪"���J?rUrR�Z�A�<�� 1��Dα�D}4	�(e��L��z�u����cs�0��-.�lDu��:��w�W
��Z4��T�� U�k����xs''Pf������gX�$��]D�<�K���Vl�P_,@�mK���\�0Z��#{ �Cd�9l���S�g>�e�9�X�C�Y�6@��nYd�"�2��NO9R��o�쬿f��%�^A�sت.�A��/��m�MU�uu/=�y��tku��PRPi%YJY\���_�ȷ�![Ȥ/6�8}Je8T�@o�`�*�'�q����|3"�j�-`���Z�j�]�2Qw��nǲ���+ Zv�g���@� �ur ��IX���C�F��x��M2qT?���`��S�F�!��r�����jҾ)Z�뜏+�kv'�D�!Fٗ�ڗ#xM q��%ܐVQ��O%����K05h揊a��PQ��߉�T��{͸��NL{�MM$K��pZ�zc�Fϖ��@�uYATŵ���>H�%:�Ȯ��ch�_�0I`���յ�I��mF]�q�!�d���R��iM�.J����(5����{�m�E%�{W�����w�L �E��vs��N�ߦ��l{q��o`9kӰ�eN�<G�_����G���� ���Gc�aIq�S���UaSP��q�h���L�
��Q[k� �?,)/�������&K��t �� ��y"�|��@_B��uu{T���4H0�i�9,�<W��w�_������� �9[\��bDt��o ��_j7��{�*�1d��X��oXx/�k�t��'6z���s���ck�[����@��,��a�J�AMTFw'ݬ�O�'���9k5�c�*�05�|��H(U�	!�,�o�ھ���_���E�
�+Nk?�p���b��HT�M���*��~ -_@�U�A0���O?�mc���ڐ����:�0���A���#}FW ��3B��6���refAR�:]��L�4N�{�m��NՔ�S���=������x��dz�!n�����5tg}�!���b/Xf��*�l�]�!b�����s�كq����\ܒ7���GB�5��x�Q���S_������-/���@|P�f4*�m
��)��j�k7��h� ����Nͩ/wR+	�F�a����~M�_�V���� �>�,-��l�Sk���;��HY��ܳxڃ��]"�����+�mv_���U�T"�� ��y.֚zh�	���z�mzj�a ����&����Y�k�xQA������Y�Y����A�W�\a����� ��dr�4���zU�bNe�˧�M�>�+�`�vzU�PJ� ���z��pl���& �y�Cj�BZ}^���:s q�:��Ζ��蛄�h�q�RЗ^�	G�i�Olr�Ag��i�}��@u����V��7�� �+�so��7c�Ά����Ɩ[7�sFs�󹦭�-7eH����K�;u�i���Ǯ5��/\�����m=�#�A��@�L�[���A?9H~���J�v����)�*5�3������*�=f�qEbq�t����N�p+KH������:»�i��������3�6��Ⱦ7{V�?���B"���Mt2[A&��J�Qm�_z���EY�e7٤��#���\B��:&o���-Ӟ�K0��4��	����|a����n�t��=�܀�
|��^��9���Z��Ux[�^Er����m���I�.�����A^ ܎B浟\Z�&���a���EO?���z\Q@��t�/+:�'�i�cQOa[;�ޟU�g�r:	���@������>�!�ϔ�����҄�q�ޙNR,�eVDV��~�|_�Z��ԲUR�z�v���M�uD�&h0Q�z��u��h����<t� ���	�|9<]u�;]ޠ��e)�d@_-sr��w����T1�t�V����e"=��/�U7�{!�% �d����y��P�A��?��.�ʟO4����ȳ�v��O\ʭJ�b�$Y�b��#�޸�`�+��]|�@O:Yؽ{+���x%�b�ͯ�
,��Q;�Y6�?Ы+ˬ'+�Va�wԋB��O�����r��(C��>���&hJ�ben��'�s?~�`���K�l�mvO�vz����]"�[����'���>y ������p� �y�B�����`�G�!zUJ�o�i��$�Mܣ��`���poOF���M��Vc��4RCrC�5�Cr��4�8����8?�ǘiվߵ��*����?.���:�`��F|C�wo�>|�(��ߺ�S���b��U>Q������5��-���;��3LI��;)��7k��v�R$��dM��"j���f��VT�V��Sy��lH��ҽ��S��oiI+��p��rE5�+�XN��Z�������x~IOS�l����J�tI�鲽�~�Go�&) �W�zm�^�<ր�����Q��-�E~spZU�@T���Ȏ!3�}�Jc�H*�<o��T�2+4(�����aJ�������&��V��:C�+�����U���oA��� ���e�.#���g�zf6��U}_�0�3$p`���{�st�`�؋�?0w����a����-�ϏO�jd�E���|�����]�lX�Չ�Il��G�ɗh+I@P�-q��9��NTO�a�Ǉ��O/���Ԉ82����霵GZ���A�`[��N�?��e6N�T���)Q:�r��C/!��bN+햆���g��h��0��[��:���S���/~M
��H;��}1vw�sv�:���ry����%���2����^��u�|0¨�nS��J}�#��<�
>�}����q΄h�@�GdP%x/J����{��b�[�9��~�b�FPr<���-��|#O�㓔<���y�`n�}�O-~3��NL�Q��Y�^�( W[#�t�A뾆t'�����kQ��Ne������w��#-� ;ˡ����l��������)Ub�KH=�a�-7�jѠ0���VP}��L�ʉ��7�0P7Zi��g�8���p�����E#��1������w��qC���Y�Lw�|d���B`+���t�X��vO�j���w�����EL�J*1�
�C�3\o�8�qX�V��*��(1��D�f����(�g4�B����I�����G��T(5��.A��/�yK1�l7��X�o��`F#1+�岺y2:zb�ͭ�iC
]�'�����8��솧��k^f�b�_���/��vm���7>>�:Lg@�L'����C�dkF������7���e�>�'�3�"
��X���A<5�&�����d�� ��?�=P���"��Ff�?jw�I1���ub���� ���n��Y��ҍ�H�4�x1O���]�Y�N���D��~�\�<|j�ܿH�ߓD 0���~��y-z�G�_���O��SW�R�^���m����'�>�ˈ^�9:�k����ubQ��w���۩f�)�R��p�[߀��t	�hNY��?�{��AXn�5��,��o��
QJM'�R.��Q�<a���}�X����7�s��>L�����~����[nO�0���w��m��U��E�//b�I7-S�HRˋ�-�-�p�'Ol,l���������7�j�?Z8.���*?+tb�O�?ƪ�(��UՉ*��z"kn�(�-X��z���J�b�����`9#�r�bW�H-O�{~�y���4��ZC����*Wdåu�z�LЅ�6068�J�g(�.�cz�k��Bxcrq�B�����^�}hP�N�K�����G�9J\��Xa׵�n��|}�!����W���!_s�Q��<���1�5e����&^�A2��J�� �K[�8�hl���1�0�W��	��F�j�p3�V� �k�0��n�D� ��8���<�Q�uG;�H���B�wm���P��w]��箿���kV�wkӊi���}�����mp�V����_/=�17���i���et��\�w2�{�XXίy�d���H���\[�R��wɼ��{+�<֖����\jj�{}�k�c�*6��=�Q���!>�@�Q�L%�`>�3�ݥb݋��d��y�ӟ��A���ug��P�wSʀ|��y�sN�	����i�0��Еc�u�(�j��k��|�\�ht����T{8(m�Ԕ�p���v�Z҂@��������G�h�s�Ӣ���Ǐss���3�������Y�܌sv�d���S�q.�a���TTjn'�V���)U*���a������4b�R�%5��;�up����w����z�"$kl��`o�-q�Z�Be�_k��m�<V*�ZW��0u7�����P@9�T<�Q��v��7�ǘ̕��7,G/}��gvWj�>Xޙ�5�3��7�{zp��t���罿77�||�|����ء�0��F#���E��5
ލ�2�ܣ��_1{_��qrQ���S_Ť,�_��ݟ�j2�(�o0���鬠�~w}�a<%Zo��s�qk���.��==������4�E�pr�|"]I������C��� �+��Y�j|9��
�L���^�}���O(*qP���Y}+suR�R���G��Ix���,t�o��C[�����0���W����Q������yY;n�9��h��� ��DG������}, З{���$Ew��8�R@��=$�
)�������IGO��I�߶:�\n{�{A���^��bt]R��$:9^��R�ҵd6��x�Ƌ�Ea����n6\�~m;a� �0����=q��)fp!�r�ӥ�_��q|�r>oa��MGl%��ٹ�@�j��J��!�}P~,[X�D��5�-e�dY��Yz�h��J$��n�o#.���A���DU��8Txy/ 5� ����n2�lZk�!���yC�}]G����N���͔�y�ڎō�T��/�c��3\�"
��V�=Y �:c�#x��������؎eoG�ݙ������_����zme��Ѵ�Ԩ����d�����@Gg@8�:N��ᶝ�0�w���E���}!r�%� ?�L`�`��_���v����:Y}w/c��@��tB�L<���	��)9۹�U�|�N�+s0���24b�:ܭ;tJn����=(��y��Eq��l6�N�yYyE}S5�l�c�LKO����{U#�ijU-*0q��&��L	�g���(�,� �	J����ӌ��,C��WM;��
��?�%�M���o��P���F$��-ぽ�վ5�����	ST�x���'x��J������c�݃�)���
�ϗ���)ɴ�u_9z��-�]�М\�+�E���Q0���nB3[�4����`�������f�����kv^q�T߲g��>���2�����j�=���Q���`~-�2�؄�=�n�11N��
7,k6?qn�/"��N�3�����p��`�K4�^qE�q�v2�68�9���t0�l`�����x�쓼�M�g�rF�4����� q2_2dPF��w�~�ʬ܏��/k1�=q�|����������8W�j�K�U�h��a`ŋA���y���S����x�r㶗���O[��8��}�_�ǿ��df�7M��qQ����
��&����"*���@u�H�(�O�XGu�����C=��p�}�V^ۭ �e.��4tI5�CXl]����f�/kq���{-n�*7��L{(i�J'�L7�	�����/u��C�y�#�ŭ>|l��n�Y�ڥ�w��2�'1WK�4Al79�i�Ѐv�zF���?�ɵVx���4x�y���)y?����y�X�.�c7�o���;9a�[Ub�~���Ep��Z0��K�D6cP�J�V� )eb7Kr���\�˾��_�?5K�&���3���#[���b'���#���&���y�&>���u`z�IJ�Z�����9Dc��v�(V���C�0�^�닌��%���TA�O����H(o�#��=��\��% &uW� �v�Ϳ�A��{()�|A�7��u2�ݾ���Q�9F<����jxȏ���_q��|�·�����΀:�l,�5�ޮ�.�_MZ:!#?�ċ\���Də���qC�d���d��bH�J�^�1������bO�#�h�:��I��G�sͺCC�4G7�=aHk��+'����c�p]�!�aM����.��-%�j��^9$5E�zY_��q�݅7kx�ᦫ�I�Ut�T�G����&����3��V�c9�O��U�*��.�/�ŷ:�?�w �ц�b˸�3�A�\2�/#N����Kf�u�<Y�1g�O��f���,HE�����+&_8��m7ڵ뫊k1�Pz����ĬKzl��MN�/qjI��{��6���s5C�(XfZ����~Ҭkra���['�iN�����ŏ�kza�&�; �E��Jς�?��V�!zX��o��)��|��k39G��lY���b�[�&N[[�^�ʈ�����x���[2������d;�.Ӑ�ӭ������i�����Q*%�жt��G���2
��}U�k��΍�T��r�k�]�by�ɞq�>f�H�~���W܉���O@�R蹨%2M>��41H�Ө=Fb>L��x$R��Bf*��V�������9�Wq��$�5����DDPF2��$�����P-�3�71e�P�^!�H�����ݣ����o�mmgdT�Ϲ�t�E`� �&m���H���@[$�л�K&���5����_�g�o����S��6����\1���8��⑲l8X��k����4J��8�h��@g�� �V���&M1�hqRPZ<Vv�)w7��+��ig��sҴ��'
��0�H����C����~���D�ϡW^�1W� 4�B��k$��,��U�q�3?9J�:�>��υs�|���?��HN�
5��f���B���*�!c�("����C;	aJ��zZ���l�3�(lCcgk��캛
�	��+Z�.�K��3���SUWě!��pQ���s	*婝�_@rЙ����OC�?vĄ S>�<���kx&b��P�ƥ���u�`}�?��Q�b���	K��Q����/)�_�� �.u��2x��뵲}�Q���,aq���y)��C@�fy_��o�?Y��1��ɄTq�q� L����(�\^}��������s�k����Y�;�\�ѻ�629�Y�3L�?�l;m���ͽ1�;pE��Q���E��-[������c��=���v0{ZU,#���rP���ҟzu�ֿxM�+�p�}��?�R�}�#6�l$H>��;��}�\;��O�&�[Ȭ�9̸I��DÅ��>v���=�		P6F�E�'	�7���A�yǵ�e�]�,]h8��c��լ=[�q������傳U7�'��-�>�h�=]�RۺLү�Qh���n��J �����������l�(sIT;����N�q�q>}��>��7H@���{�%���"s��$�{	�w0�+~�p۹�� �MT���y�)Z�Iۚ�z44�������%J�u��Q>�j�y�+4cN�P��L�I^3�,�ad���L��z:k'�Ή[;
ۧ/�aGf�eϡ�A�]�k��@�Z�!c"�o}<\��bI����+�b|p�Ch�ұ
��v��J��AZb����"���#(}mE�z��r�6���[[wM��`��@�2�)%������������]��S�bL�P�X�M	\���̅9z�q7���lܠ�d6�'������q��������2O."�]Iv�ÖJp�fc^�5,�`����������A�R�zE/j��S�X*�:82n�߰�����ĺ��¶�ǩbQMP
�QW>L-��W���o:�OD-`<e��i�}[Υ� �\vb�k��enk$Z+�y$��R�FJ�WW�ǻ�=�C����q6'v���������f$�䉯����iU���u�齫���O�W�������l"u�4�߈ �ڈg��$�I���;�+����(q/J1B9��,[Sk���*���/Z�T�	 "�@Cy��1��g܍S!@�˾M<�#��V�N�0���K珕��͝���Z?4�h�������=h�:����B�<��;gQ�HO#l8B�h���f��3��GVf��4P]~�m�4��a�o��[!�5,�;�ʐ�yS�Q�5��H�<�}�!RC@�4#Eԓ�l��jab�u�����a�+]�}QD��ڝ� N����u��3��:L>�����X��hH�7&��{�=	��{�z���k�r6�l{]eN��w'g�r� �����DlRLT����7ʫ�+�K� �����N�?��5�3]�{>��z>(��(�(����k(�_gf'`e�ei�	�V��I�N������ބ�@�����ce���eN�#��~^��k�P,��}���� �ǽ���K'�"Y��u&
Cd}�w�iP�ڕn�)졟�5D��tׁ�:��0��|lQ���\.Ɂ��q�WX�h��	�+~E�?�XR�.{�g-V+K��q�QL��`����ꛤ=�A)d$� qȡ��" 0=��?��������m0��xSGR�$z�����[�Lp�kw���ӗ:ݡ���n;�;G����K����N��%��~#����v���91��x�5+���7�^�s�e�<^�M���%�$Nx�g����<*��~�^EAtep���($>�Ȁ)��T)��\��a+��!��^/�W`j�1���g!?z�%����^Wn5�x�L�|L2�����G���n���ݒ�yY�Ha�R��q��u<��a̕�5#�~'�6�_u��t_ԯB'[�Jf���h4>6`�?�x-�g��w�Z��Ш6��
������f��vIsH�V�N�F#�ɺ#Ėk_jX��/0����z����f4���g|�!��g+�'-�a�vE��3�T��c�J�+F������RPpÎ�ǆzk�':���˿����GQ��-t=i�����.?�8����&R�a"�*�e�_�s{��w�(�]E�[_ߞ�g����5�v>l�-z�[�cޠ��o(��˧Y!������(�6=гX1�����x�0\"�Sg[k,����CRM���������I����(4`gË�n�����5]�1�V�����gJ2Q�=��#��]��K�^�`�  Ɵ�N�n������Dؖ��D�Z��;�,��kA�gY���iŘv��;Ǧ���s}�V���nw���Ѝx�y����Z�h�c��o�M� 1YrU8�/��E>9�(��s󝸹=n�hNh`�uT�K��e�Z�Ybc�˪�C�;��8��9&T3��+g���!<T�6�j���JN�	Hx=�#����o �n'	7Q̚ݱT���$-w��^����mg��K��OT��%k8��aJst�5ϑ�ԲZά@q����Y�2?U��[�8���4 ��z�3�p��Ah䡞�{
;4
ޯ��*C��k���4����c�]Z��X_E����;pE㵡������:�������?�#�ѯ�J��w:��#C������#E���42�(p`�����j5���^��B�vxw,!�|4.f��R�޿�o�&���O�&[��3ʢh˩S��@��m����a��~^��fD��գ��rݭ������/*���OR��+����2Pmb��"��"B~H{��bm$���h���fJش�Z�RL&���p��6�S�?)^n?9��Vz�n�hWdZz�- &�e��2s�-B�TDa�ReYA�x���B6�|%��������YE��jk��O�����$�`~\��4�b���`	�R�A��ڕV�}�77�,�k��`R�Ϯ�q�a��0�%(d_�w��s�1��`�$E����qnt��I���Kq��u�#Զд��Ud�����zK\�}�"�Y3V�hOE����.��̆�+4������=n�m�zr��$y�"�D�a�9w������;i~� t�����ΏM�u�_jEu���5��-��,�F���eSU�$���[	Eiׄ���-GkU�{`�v��B%Q5�Yu
d�(����B[[����w��I#T��b��C-,K�00;��&��:��R}��[���#�v$ �,���`ђ�E�n�jԲ�=lY�ٸ/vv�6
�a��cg��r�ֻ��O�FE�K�~]��,oWK/x����6�:�(���͈�m#]�2cj�^����.Zo�pAੌ�)2F�mÍ�-x�� �vi/�l縛l/����C�W@5��������R�!!*�J
#��H�(!��J���Q" �G�!���L��ϣ���9���x��]�~v��?�������\��Tj鈨�g���1�s�4!�$��Tɪ1z�.��NL2���N�*=o�`��N^����W��z�\����k��uꜩ�����[�nk����M�d�p��7��@��"6�PI����N{|�u��\��	NG!ӆ4�߇4���y:eb��q���r�8fڻ�%��|�x`@cK��n����KX�7M�T�AD�,��P��	�0�N��Lq�`
0�$�Δ�gԹ��y���Ip0&��b������y=麤�T�>ǙB�;��5wd�׺�b����)7�˶ۛ�m��	ƣ�����^t�m�`L� �v<ꭺ�s��}]���3�����bD:��[�S]�ܵO�)Hѵ������{B��H����B��}#]�fiB/�%'K��}��D���M�s�����ࣳ�L�l=��� �=���(�:7�Z�����>#}OPdx��.GO�&��"���W/@'\����4'` �b��Jms#S�
[i���4��HM׾�K�:�<%�YYƶ��K��ii��<iPa�a7W3(�@�ƴ��0�s�h��"��5ϜA��8͡=66Ei�w��Xq&<~,m��G4�9��cV`�)[��ޜ&�3��Ѡ��BQ�d͡�|n�b�B5,��[F���ш���eە�yh'-���}(�4f=l{��!�R�[m��a��ic��J-㽕�`��R�f^�31~d|�)��ו�"Phc��}�����Փԭ�JΕp�7v�8ڻخ�t��5Ui�=�i<<��ڹK3^��l��� �v �Zvf1��5��y��T��&h�?����FY�EͫVc�S��ce����M�݉jme�%�q��^o6�o�,0�B��M*��i����o�yzw�`�̊�����B�]�gV	��D�g;�w	NL�'�V>�_bj��xa�����jB%D��&�����V�@'`��F]WHtLӓD����{��/�=\I�]��_��X��i�Eii[*��m͍����o%r뱧�R�'W��|n��d�A���J��&�>��-e���hr�=�[g\=��!Ot�њ@���D.[+���

�=�A��|�������J��AQp5+]�{�l�����c)�h��(9|�tY�J	\fڍ��C�p;�.6�Ą�?�fK`���5�3���{FOG'�:�hm�K�,))t�k���u�s�=H���ۄ�#/|בn4��۶6����8��V�^����L%e��o�T���Kno1,�����6�uE�g6�w,3�\b麌�k3�&��{����m�Z��F�͑���ϥ����S�2�˚P>>��&f�8I���I���B�)��k��f}��Y>#*
��e��a�;�{4xyEƝ��}�C���zQ�y�4H����aa^�j��Z:#����U$���N��{��n�YFD9�W;_�v��ڟ8u�U�f\E-�?/&r�-�z�~B�[~����AW�VZ?,-v=@�õ����s����{0���Qf.�;��t�k��`h��v��<��Q���*�>�,��G$�U����f�>y
�m��H��S�z����<e����u�
�� ��5�C�tf0��z�IX����g?=�bX�39@��zl.�+f�x���$gp._i�iUrɀ�`�2u�'�1�	��H�A�>�>q k�xw��?\�^�΍�����D���i�5T:��#+���E��,�z��o�7�Э�47��+=�Y���N�.�ۧ#�U�^�U���VL�*�K>J�g.�%���Bġ�#���٭����A�ū��D��v{8�Ҹ��r;�zPjmP�7DL��rKtV�_#߂g#sl��C� T��n��d�����F�S�$�A�	�fܢ�-��p�uZe�]�{�k���Y����z@�X��鳣�%�)!?�3\�dBǩ�#��uX&*$L绰��fG^L��)>�|�i_�
�1���h��T���I���b�ݶ�
�
J,�	Qf���}mX6��U����6i���̢X#ޞ6�m"M��eI�?��%8�M��O>�s�?�����,䲴�(�����|�m���o�
+��#d�elg�+���O�ܥ�
R�_l�SŌ�J\=�BYgF�q���p��������:�/����m;E���([l���$se��� ���xN��)O�R�SO�"���2u�;7d= �>*/�N�5dKܽ7�٣ڗ�+"k�}F���9�c������T|_����E���[hH�iAd���YT�
���-�<�V��cޅ�aߚ��P���{g������Ω��y;Z������A;FtJ�����M��CQ@j��(A��ׇ�e��Z���]bhpX����>[@�ؠ�E**�6^g�lĵJ	��5B	�.�o�\�Y�n)y����a���\t߆&��pjx�ﾰ)�ҹ����<�:˙��J�ܨVu>u� a?T��kk\&1����
��姑g����]_�@H�SlGtun��h��9�5F[����c�@{V�g�%��r�����=�O�{ڲ�!���MǙ�u���E��5�3:�]Z�5H�$ҏtҟ�r5kO[6�tKuK�:\4Kj\�ԩ�.����C�.�:ń	ϧ2z�fAM���E^�.�(��O�}8�9�������S�L�2(�#ص���O��s���Z�AJ\3vI�)2��H�2�sPb�/dB`��9UX�s��O�n�N_����E����dw�w�N4��ҹ�4�R���:�H�����e.�3�k�vԇ��ڱ?L�Z�@jp�F�0�A94��U�V�"`S��5T�\D���:-�08���f�#S���~K���#���u��o�,硢�V1�o�4iL X�Ta��}u�r�a̡F�کZ�J��a�γ��I d�И��o\gLl�����9揎�t~�Gn�>Ѡ5�>��Jl����2���s�B�if�'�W�$��*s⧂B�P<�$HfWT|�u��%�Exٔ�|���C֑_/���5G����:	5� ��L���9�䤎#���?rV!4� ��v��GP�F�Y�H����mC'xl��W_4��o����X���X���F�
/Y�}���
8��7_��W��G%��}h��D7�^�\B�'�\A��W|ۯe������,�y���"�њ썝ȇ���[,r}�Ӷ�D/e(��A�U���c�;W/�[m�<�G9��(���6�t�OR�h����߆
�7ذM0IxΩ�Q줸]�z���X�.����(�c�Aw�iD��'�������V�%��s,��r��U�*&�3u���iZ���p��֋Mw/,��j�}��e�e%��C5=�c+N*;��&L�WU��]~�Y�R�ι���۞�귋Q�)C'��L��!j�N<��������nG��A���n/�����"ڢ�F-��ٻ���.U�k�;�4�'��p����ю9�N>�A�{���R)��v����TI�?�2$�i�)~��7�=4 �9�w���#I�-o�����j�ޙ1��hE[�xaUTm��i����T�Z.��.�*[�!�.�O��Дs��Sk;����{�
�?j;^܆�nj�=�&�ǉI������695����� z"&٨��
��0u��dB�t]I�khw8����G��Q�wMK\�l8&؂ �5V�47�3��.3#Bp&E�Y�Gӧm��v~��
A�	��D��� �!ߞ�W[�����B�,��4���'��v��o͊��5�i��4�
�PgS���vU/ �1��p�lf6Ux�W5�U�b�k��F`?����&rrȈ��-4f�u�&�	��V:��D�h�dKΊ?�V_|ڋ�;ŻA��C{)����^y
��=5w����M�o����b@����^��vt��(��qK:#���͉ 9�y���:�g�0h���$6�K�9�'�v[���r����Wr܃��Y(�-�IA��c���ah/��X~����K��k<�n�i,��ښuT�����IU~j']�e�����񎾓>�HV�]TG-yU�ߘI��;��+ٚ�i��v�5�[�=�t�"�DB/49痔j=Y�9H%I�]%l/��DN��t)8u��u
P�w�����*I&�#!)Qp<�$�vi����G����]����0Ѳ#�g&z[��\ȍ"�Y����+��X��d�1���A�s���o����ãrnޓ�R�%334�L6e!k�a��F�r�P� +��Oc��w��sn�W�J/f�"Њ���<a����.g7���*�=�=���6%#R]� wG;����O�[��8ҏq��}cP	�?;���(e16ψ�v�T/�<"j�vq����6=�ڤ�	W� 8�����w'��wdPׁ������M�{7_k���u<���>�ʲ&/I�s�aa=�
]��V���r�)`�a�/UR��z/Ȱ@�>	?`�0G#�Q�.�#��۾ul%��Z�^Y�e�0�[�(�Ro#���י?6#/�#����v���$���e��X?C�*ٌ�@#K���U��&��,g8��I�u_��LL��,~
ƏI}l��g3����K�g2��P�[�hj[y��x��x�K]_e��������T�x`�����k|b�!�~��D�2�tb��Nq<v��f��wq�����1��o-,��w�����^���t���I�@av����Z�e	^����vM�C;��A�-������}̤����$CP���ϩ~N�5���$E�9(�>�qе3��,js�9	?�Q��^�� ��'��nO'Ӏ��Z��m89�Sv���W���2�l-C��Oj�!W���^�י�|h���+��+��tpN��k�IG��F?�Y�d�����QV\�JJ2�Vl�5��)>�w�������##�������Ș�	����?�;�-����|ը�ZS6����'Э�ܱ�[�r�{�{<�-0D��i��i�oS �M�� 
�t���������o�A&�*��vĽ{}V�����M �S��:�$?�e�R �)��]8Ѩ��1�k�m���*/XA�H�b[�\��x~�Ap-�]�Qv�.��_�9�(�h�NV%0$�,�m@����R~�ըMY`�V@ƪں\��@�
�ƪ����s~):h1��w�-��W���r��זzuߠ��gJH�	9j�+��)�N1 3f2f�m�w���.�&�
q\-��.��S,�qaq�g
@B�ʾp*�|���kpj�Ҽ����8M���e��G���w{��;[Ok�;(��V��$���(*O�3�M��#q�_��P�C�p��7�MR��&2&�W�Pn���隈��o���'/�t	�|�hJw�yZ��4Sf���F�pQY��c��*$妰K��6_�9u�����"���L7�*�/i�M2����y�ĘTL��ܠkP8Zc��d��
c��C�DI���l���6H�ˡ/�jVSKb���x�R&iձsy�j\��B�����{�}X������K�@R���C��g����;�}G�fc�CU�/[W���I3�C�:'D��_D���B��������Bi�N�i��I�V)�{�G��D�v�(����RoSp����Τqp�rp�;>�SL!��3��)��b1��ͷ���bw%I{t+����;p��������'�������fb�6�{p�:r�0�ĺ��3I�k�{a �Dm�� ��6k��_"և
^a�u'
�l�(���3`s�P����_�U?yf9�]X>�e%�#c��Ú�2�'���"ۨ��j��i��;�;͞&�s�R��k:��v�[�9��h��kgI��VBNd!��Nw�Ω�	���Z���yr�BL�ȹ�4(ǵ�ݼx���__6ɿ����;�C�o���U��O}�4[�%�l�Ae�z���IžT��'t�>g'磷v��}MczL<��c�`��u!��a���=M���cQ�m]% ò�f˅EHe���?d��hX����Wڂ����y5]� Hd�,j�����\��j���՞�g���p.��Š�=��]�?����?:��^&4H���w�d�Q�5�D��E�l��7 ��`���@��x�<'{.����A�޾b̬C���q�N�G�_�X�a�݀0���]�G�V}���骦���J7�t�yul$JU���/������a�I�D�-�پ�,��R4�m%�Ɠ�d�
��K����Z�A/��J}����8���=�����H�~��p�C��}���q�n"���g��M����]���aҐBt^�k ��P�����P�޷4��sR�����%��y��B����"�=,��q���f֚5(L���\�FM�*��Y􃶫Hl|n�}�;�Ee�.���w����{LU�� *��E�CS� ����B����өH�5" �͉�]|����@�n"r=S�D��'9f��Ѯ���N��E ����,l8���5,T�0L�Ӻ������ǈ
�$j��VZv�)� bv����������Z�w������kc�;�oYK�o�l�Ԣ����#]�����{,���(ΌcMs,y��$��B;��+Kj�9=1k ��{�­��ݥݫ΀�+ۊ�����tO	����i�#;K��!�k��4�d�Rg�+���K���z;�*��9:���r��@������d)��;C�W���M�s�9b́�FL���t+@'@�Bɬ�)748X��-C��`�H)����x�麀a;;��ӂE��/l�J�Z�F
J���^�^2T\��O�op��7�s�LR�s����? �7��-�e����h�Z��ᩔ;��q>ϘxVZZ|\�}}M�a�j��r���FT��۷� +�g�_��^Eõ�ݡ���<c��?�=��q��R����NOȅo�ř��?������?��K�p�#n�C��WpAяO��Xw��>t?�ņ���1�	�ť�K+{A�En^غ}Q?�޽�E�=�R5t�P�oG��7���?a�l�+ќ�� ,9:�=���w��L"D���h+��h8!�s�t&�;Zc�7�^�����C�GMp�D���z=�2D�9�J�tw�(m~���57�5���㌭�^�wC��˗*nx�}J8)-E`B!�Y(^�ƙ�l��l��Eҭ�V��n�x?�q�"�'ZJ��1��FLk�fD�<C�@�D�����?�4��h�LT^�5�BD��fq�s������@+�c�����b� "j�[aB�=���?��p�d��T��@ڢ�[ozғߊQ�o9zk:�nl��H���їZ�����-c$�ҿ�N�����'A#������4l
A㾎(@�1�ԈA�P1�2A�_���>��(�|u�'m����4Hb�n���L�����k�g�&d��O�j���z���'i������=8��#.u���1�z#�	��c�ȣ�5�SӞ�H��k �h�S��G�p�Y,�U賹 L��=]~��պ�5����"���ޛ߁ic���lLy�ƱXT5ҞF�BT ���5%��ۄ�8
VxAO5�f��[�����~���"������&�����y��1~�	,���@Z�!-Qf_g@�|F �7�l��y�qt{�<g3H���_�R:��65��+���T��[�Z��]�I<��+�D��㢗�6ب6� ���Nt�,xOS �.������b
/I��S��l�M���&��r�#�/���9�Xߋ�e|+P@>�;�Dc+Ep��1J5$�m� ���H_���OK�Z,�/p��B�\h ��Vh���LpXϫ!p���Rpw�
1�e����5k�dp^�3�gn[��n3uB�M��O����<%�1d���G���;��K#D�;R�~�~�/�34U �׊q�iX!L�A� H()�L+�_
/���~��cď�
�ӓ �O��e5�Q���ɻ{��c�����A�E�_�>����U'(���oQ�:3,�1�o��|t6窻�`�y��_���Z�6ʂe��}�n˘�>�5Ď|!����ai�hs���W��O���g� �-�c�����S�㶑'���
(��`��M(����%I֍t�|���C��3��Yw��~������5�l���S�'���|+��{'���nc��$����ce�G'�S����5�����G'o���v�����/Z��� �|��7�v���~3�B���c|f|�Q(1qB�q':��P�5�>G_��[�67Y������x�`7鳹FX��5']���m�Iʁy�Y��t��HW��*��!��?F�������dn`��c�T܀� P��0�����4b�M	O��H����+�ֿT�>i�Ox���ocl��>���o9諟�o�P�Q���2��V�6�������4ʷ��gh�|���&%f��{3�k�qd�oP��6H^��r7s��*ʅJ��}��{�s��y�.���?Q�#.����/���*_l�Ecjh���#B����@y\y���{���ci�ǋC��PU0Ah�ԯQ
��'a)8؋;�;o "��ؐlͦO.� �
è�mi� 竫Љ7)�^R�S�$�P�J��3�2�Ej�?v�q�����P��N.f'��n）��x`�������	���~hj-�|G]�c�/�˰|��.�Ogk �uь����US���~m:��hY�ђ_��z�j��a�l���X5�Z!��yw(��V������U��NS�>0&� ���ٗ=
��QR��!�>��-)6��MVU �j��jdf�� +�U����Yȳ<r��1S���{�-���\5 "�,B�g�HA��N�P�0b�x!��.;}�`A� c��hqy�t�Ե�@&�s���Ė���y(@�*4����|v�����>�6����0�
��������ar
iw�.{��G1��l8w�O�yd+���F�P ޑ�Mr�'��:��Q ޝ��h,���  s�q՞{?�9R"o�.mI?�+�T�����9����S���8F͟�S��G�\��F~P��)^��DD_�
��0\��������Y�Z�n\�R(N*։�Ϧ���gO�N8б02	�3tt1,�E��09��>! |�����W���&c��Y0��A&�#����#�������������{)�%k�=[L
�c::��B�or�1U�7�#i�ב����*P�		N�n��d�Ld�@ܾ֢���+���>b5��Q��ؤ�.P�<�����/��jhe8���ѫ�?�&d����I��}ۯ���������YЫ�me�e�.�`����-k���ʨ�it[_��+��l4��c�xi�O&�$���!�G�ǐA�W]��k�Cq���Fm�\��PRK� ��@uȟI�/�����2ЋRL��g�uL�6�H5�ʵ$�+��B�0���g0�k���l��?��U����1�1T�Ւ��7���\����9ɠ&�v�,#|Ye�u�,9����$��9)��"����6+tX��~ΞLI])Lf��S�`�xw��67�D��8�'�����MZ��/��)������V�S;E
����_k�	� �o&����x�v<\%~�uP����)�v'� ���85 ؕY�� PU����Gǖ)v��Q��1�&'��V�Ś'qi|��c���"��_~BE�0��.��t?����|��k�M8�@�Q~�M�9�ec�B��ꏩo1�t/C(nQ��tYb<"�fMד��z�>Wa�|�0�����/�6�ܙ��q�X�S��B1ǩg8N�(���;+��@�͎�W�����|pAǦ�$��i�-��0=tb1����d4ڏdL�B�#�����2�����]��R�3LPʗ�8���6�}����[\�T����e#�<�f�|�>'����'V�Ɋa-kO��2�������������eS�;��٨�1&N�#��3�����O�j��-Z퀬<�ڶ,#~��i���iJ?��8�1B�gvB���WIjM�79EU�X"���ɔ��ɮ�B��v��\�
��E�����nv�x� �TVey�W� 	�w�dƁ���
�^,���1����p05�Jپ58=�O�nHJ(��{����j�7���|����f4��Z�y�Lʃc�h�T��#�V,�+�!3�qsÕ�@>�M0�����~ћ�D�M��o5�s<8k [}9���م��~��I�>��ŉ�9����h�b/�@(���ʫ�8�`����r�;a�L��}Y !J�Q4	ԙwd�c�[0L�A�F�j���H��ey��l���y	���扉�U N�m��g V���9W?�oNτG)1`�zr�[Y5q3Kw��1�P�8���U�;iz7���-��4p��n�D��OQ��ϓ�:��L��Yple^;�Jhb� H����,�K��n-�j�� ��g�@^Y$��ZǞb�_���W<�b��2� h}��r��q���e<��AU7�}�T��m�ݵ�^�)2ղ��RM6�I4���W}��cu�s�wv�F=�F9r&9�OG�Rr�J��j`���6@0��)$2����5@>~�Y�V®��g\d�O�Z�A�I�B�uT�A}p*�\Գ~,��m��������Eh^�zÿ[U@Ywq��'r�@P	
�U@�m��O-��KH)d��"��$3)6Wn�2��v��}!��E�V$�@Y����hKrL�܄��a��گ�Rf�M�I�TxK��kY��n �*���b���0<�G�� �*��ͥ�}���N�7W�J4�sh����
ǃ�A��`䯅>e��*����L������r@x��X
�D�d%����[�2XL�7hpB�m�ɰ0|�
���aIw �C2�&vVtc��l���pI��$��NN��~¬E�	���e$�h�qt#h�^���[� vM���e�ź�+�)(��j�������Ʃ���5���i$0�3#�@�wQ�`�Y{�ϯ_��N�\����%�v�-�d_�����R�&�Gj��Oo����,�7���r>1H�t�Y���g{��M�dF��N��Ԛ!ǡ�<Sx�j]�d^yK�ڧ�!�u>�� ��4|�zN����u��V�%�	��y,@��kp�r��=��Fe�H91������|�Ϲp���5Dԁ��=�&{Y�g����<9"��(
m 8,t�H&��Lދv�]��p�jl�x�\v��|2=YW�6��z��" D��:D��O��R�F���}�����&\��2T�a�8�r�҂�2X���r�.*,��}�6���4�Y]@������Z�xqw��j��G��)�-�n50���|g9�B��^7p��4ӏXk_F��MG�tU=��ߨ�S�FƠk`�.�&�߻�Q$�����YQ"�r}4:��Q`����X�DZkx�jc	 ��ό]���fɑ4�iRD���8����UZ��6�i[��w��0g��"4ݲ�D#�J-O�%�'��lϯ�̞�pUEp�ďb�-��YT�B�{
��n�㙛]d����e!p�����d�*Hn��S��?�b���G�ƛ��
�(��H��.U�����R�*>�9�I�jޅSD�WB|s.47dW����T��fUvrt��JFҙg8�g�c=����Q�Q��+B�Ŏb���tJF�}�-����ܻZӪE���o>ۛ��I1�
QU������S���6BWB@j�����`S�o�����L��Q��lx"��h2�Q�z� k�@���)OYf�o�T���M�*��jTB�B;���Do���IH�Y(�NK	�yl0�ƻ�f��w�mG�0�L?r�Գ���#�òБ���$h�E6�:f�q����4n^�ᚇ"i���i�X�Y�M����sX��fҽO�[��-D�߭���\�޴ԍN�jkʅ?��w&,+��<�fJ�U�Y�>'�7W�w+	M�Eﹺ��8kV�?"�6��շ��N�Yŧ�2�*�{��i\td���_�=Ox�&�|�A��NYZF�����`v�~�R)�-EA�Ɲ���P*�y�t�꽠^�<x7�ٌ]�{{|�)i��`���'s���+�[��ko/�y�U�7ܰ�s0�}��y�Q�����}�	��ȥ�p;��#�ר����dj��x��w���&����PxƤ���N�U�����j*e-��*�;h������p�he��i� `�����}��Ү����+�X����,�K~P�R��N��Jt�˪�[Aop�Sh��r�j� x��|l�Qߕ�+)f�S�]��-���A�߬h�je�Jfr�/��UK��$|�1��n�'��o�$7.�H�@@Ĉ�*�V�=y=���GK�w�������	��92&?��ͤ���Cp�#ٵ�Ρbk�j�:���@C܈}0�U�<큦�*G�������ҵF���\;y�D��l�>����r~�+U��lmh�B�y=/0v��S�~f)�u�ԍF�0DRY:��,#]UJ�x�?��k[�������7��xG�em9q1M�_Q!4xb�hG!`:��1�E�s	u�O ����69<������n�6�=^L���,�}7A��2! �G.��+�Ӿ�w��'L��<ü�c?�3��ՙ���&+�ˬ��&_�Ũ"#%�lXs�ۙ>X��dqhK���5�U�/i3$h���O�N�b�*�Gpl�;��z:�S�_��F-M+:�qE$����Uxu��}�8��7nwGh�������.����}��0��TE��%�	����}X����9e��Q��m���v<��3y��/<���y�?��#�gGӜ�lby�p`��z!��]h�C�_��"G����ȏ��4U=��ɰ�7E�)%����2����-;���4/�g�r�Ɇ5��va���5��
)�y��+!D/b�oMC��������@�OKI���<c����(��l�p<)�l�,�3Q�a^�=��{�f���!'fkK��n��,��X}6LӑgI:��.�@U��S��OdMHu����D�Q�Ǫ]^<^c�;jۣ�P&C��	5�k�m�u�I���a�ö��6o�|�����] m�	���:NP���7B�Uo�z�U��s}I��ۀr��O��4<4�}S{�'�]�Dw(m�g��Yl��i���$�S�87�R2�;-���H/�Zڼ%�J�e'��衒�^���͗n�|[B,t��]�
�=�?:s��>��ٕX����~ۢ�Za�՘�1H�=��J>Q�\��������S�;4W^�<�&�m������x	�C%�x*����"���d��K)׵P�<����[�3'qW��<M����RA٧������9�f|"��x}2[�1Uc�4�@O3���,7:ͮ�cӨj�f��@9�u,u�#/{�J��rtYEpA؍�y�v#�%`�i	���Nɪ�WΓ��뗝�味[��W�|���L뷖�p=C�V6f��7Ҵt�N*�s� ً���V,�;I����J��1v�2���W��`�H9IAvj1���(�w�����^�����o�1�.x��kʛ�>���t�~>��E�������΂|����n�*R��Zb0O5����K�g�z��ܤ\�ۃ�b���,��n��yw����PT}���T !���:�cc�x,OD?�H�茬��E��g����@vQ��K�2ń���{Fr���mo�YvN���xQ���E���^��� ����3��#�gsA����	X���ok������-���>zy0l�#l[l���|�CEa|�Qr��X���~��F��	�?H���x���=��z�i�$��ӎ��9�e��f�(W_�������@��G���B�\i5=���cf�tBNA�jl�:�~�cl� 1�a�o���E6��/��W�������n��{2�&>��sv�`��~t�&[*��8!2"���-�6����Vk����8�6��$���2��Fi�k�i�s|G�p�Z�	��jq��d%��}b\���iLv�pRƸ�}(]��ϻ �U��i�<I5�h��/�@ʩ�����fx�k���@�δ�F���w����x$��������(ԯ��o?t����V���[}����z����,��D�+Pkf�Ρ���f����C���%�|Hl%��	����N�m���SQ�!����(2b�<�}v����;XP6��aUs/|����7)�hw*ոDi��~G����������2@Z���B�^�m?C�a�N�G�Ntw�����Fa�����̔��Y��X�P�����g=w#u��sG���D�Moi��^�G��g/]�W6E��:h�RG��!{k-k�s�r����h�P�����Bl�*���I�q�M���M��v�â@��ǐ��@���z��F�`��!^,�u:b��ݨ�,鰕N���l��H� :u��G��	_KTZ��{�v��6�������Y���U�~�[�x�O߇��,,��J-���t7����QVtb�����K�6"?c��)j������=���F�Ϲ��ّ5�Ra���q����r?���Z:5��7�&?0��x��������|�	�:}���r��+�IQ��0.Ҟ�E�fdb`Ϟ�*k�Ў���$��89��^(�@�wծ�"+`��5-3�7��ɣ�e 7��,���Q;A�2^��b1��ۯMq��׌a��7��{��4�
otB_
�J�ğ7�3!Cvg�˃kʐ��4#�H#��%���=?�|�+����n��ҹ}����djڱ�5�}b��Yi�wlD̒�A���n��.c�iQ�}K�.n�"��ʳi������nX2����-v��f�'������Y�>k�RL�O����O��<��k�l$Gx�p�$�%I����Q�hWe�/�?��P!�9�:O6����ڟOc�O3_�W�.$JS����*��}��뤶gs�8�w���L��2�n�9oRvŠ���:�3*�Mykә��:m?���2����:��Kĉ�o�}���իz-�t����L�W!�Њ�`�"\��_?k?!v "J�����9���1qN��k<��]�ZYA�r�v҅�*�}��Ft2ts1���8X����[��F����w��D��E4�uG�,�~�I&�����ƺ� ��Q���-oO���Ԅ�
����&�r�@�2�ȶ�{ri���k��E��p���u�s����t�+QS�s�X�
tޒ����R��b���h<f��5�^�{+��RX-j�Z�su-�J�K0¦0���m>�yQ��?i;��!�����4�J��u[_��s�C�~_G�yM��
�%)��N���c̈`Yf�w�������֝��[�q�S�!1g�}�Ҽ�z��3��?;�B����iT�1-�$����D�y�f��F�F�����������Gw�W�H���i�x���Wj�9N���������S󐀭M�V��I�����ݢ�i�aQ�d12�]�M��K�D�@����^��`��csq�� -�6 �e��:-�z����� s�Z��-�X�Y=b�E-���5�++��?����Z+�)��	Wh >�y&��O�&�����J��t��T����>J��#�*� ��v��s�C�[Ֆ&t�o�;�%��vߕ�}�Č#<�(��8f��V-A��h3��_]>�wm��S1�:�+� �\��
�;�:��&fSq�b͗w�_/a���pBŌN���J���'h��˸�C�(�,�ƌܤ O�p ̽w�EO�J��K��0�}Ď/{z�%=T����}�t0Q��K�_Ͷ�� ��̤��#�k�!#o|���Q�In7v��/Ƭw�?�80�1oR�jR�q�h��,�u�}˸��7�������"s�z��� EUXOv�Q�K#�Ӟ�n� �&Q�����i�з)�yEҗ��sb��	��Fǈ!���N
���ya���6���P�8��{�Ǖ�Jx�o��3�(����[U	�`f�q��⠇��h���DpT �?m"~�9*ު/�-�ؗ�A��5��uI��%j�ݜbI|H���������6��6]`vw_e'm~���ۯ�~����l����yj�Z���aN���9}u��K({���{5C[_|�@��V�˨6�����H���:����l��P��D�z�L�?JǠ��r:�h��?�n�l�Ѝ�}'� ��F��8q� P�e�W/��%��I�'�]
�6��6�A��Ԡ-}���=�g������dԙ>KSP�G~5�s���OY��!��t8P�~m��ŧ�q#�lЀ��jڟ5oF�Ο����qq���z�u)a���To��y��)eo��N�xn���R��箖��mᆷ��x���Ta��=)׋�I���c�ӄ��O��DD��\CZn�XXi����6%�߲ap-m gZK)���5(�!�s���b_���Ъ�w�f���U$�3C/����k���(�հ{:	�7EZ���� ��<�_�S��9��&����<�!��}� ���}�X3D����d�K=Hy_C���c�_O���$3d����o�#�$5��Y5�	������5�O��`�&PS)���V�;#��ݧ���5u�K��~�=�7!�?I�m|y:�q�߭���_�����V������(�a��w�e���p��z[J�a�7Ǜ�5s�=�9�n�(�"W��J�h�?�;0�$x0Lu�R�Y��
T��� UE�i)�}��'������^:�L2�X �+�e�2�`ؘ��=u�/�i��N�ԂG��Hݬ��W������~{��҈��(*�׾���������1��T�������s��T��ޓp���2���^�?�h&hզG�7�2?y*���G��5����g�����8~��UĨ��"� 	9)���\�%��`7v��-N����(�f�؁���~S����q)����|�r{߇U��U�@:DPR�j��=H�P2C�J�H�����PC����C����<��?[��?��r��u�u�+���Z��I��x^a5d�R.R��%��m99[�.���a���a;�6p���	UUE��)�.<��`4��OS)@5�4��P�_o̩�ʥ4 �^����<���v�rX1�����53���zC��n����{sxn&��@�s
v��;Z^���j��ɺ2�K�����7�����E���F-����j$��u��	�6AY��t):����t�������RJN}��pq��?]7����|�vc>g�ťiN�O��_���Ͱ�a����RǓD���q39����y�pŔ����Q��j��d��H��K�ȏ�DSL�c���]�����C1������}?��-=^����wQ�q��ﬠ�G����2F�!*C��ZB�X$�Gײ�Mm�YfWr <k ��~亷d��any)@�U��evR��o���	�}�,,'9��R������tuK�R�w!�/�/(-����,34F���B.fW�$C�?�T�M8� 1.�
�I8{7�;��CI/ז���7-�u�ɗn��Km}�?h� BI�|��hcV5�Kqa��V=��?x2pR�Dr���=��0�иjL����Y������ň�T; ��6�ƿ��
\P��3
�++�cu}��x�7bQ1[@�-lU`��o��'�:����+��v-��	;���'m�Z��~S���16ߺW�*;,<�k�˱�$������~?s��M�Gw���R����rt�.�Ykv좪�9���t :�������4��^�&
�bt���|���b8����kH���K��Q�9��<�;�i�<t�#.���L�pT'��x�Ԯj�9J������!��#@=WjqsR�36ˡ�[��QߣU���4C�OK���ҷ�_0����DØ
bX�0�͗���S�}9��6m8%}rm��(�<���dm�WX���Ƒ1A�Z^�4��}�̤�� &���UI��E�D~����n�;ڴ���)�0��m3�`�ۜ��D��R�(��uuX�^�4Ɲ�����Z~��I�m��z[e��ӽCt*N��-S]�Ṣw�ؕ=B��f�����*�c���e��7bv�\���>�ڌ�2��
za:���o^�����;U1�8o�bnCJ��j�0���������3��W��*D(z�c��h����n�d+"���1�y���M�'��]��ge�9�9�8���>3�q���B��6o^�y��^in)�����r�>M�bb�� D�KNK��;j�6��������^�h��Tl3ˋ��9��� x��`��f����*5pQi5��ќ�������>��S}nG[���$�:���k z? �?�L�tP%\��jY=���],�t�c~ߢ��sQħM}C�Uj��U��@c9(�4�5�9��ҳ�t���`�^ˌ^r��ǟ%��_|�6��+��{/���p栱��̐���SCaA�F܌��>�Y�L��?.��ќY?��Y4iq�b-�'m�򭬱���^���s��n����Z�r�\V�XF9�<jh�C� *ol���]�WR�u��(Jw77���G����~0ǓLe��v��(s,����-��ƘYi�D�ѡ�B��jox��? ���y����4d��{��(��i��Ծ��$�r��1�'�?}���p�JF,�����r�d8���[$�~W�̑gI�3�|{�̗0��~�������G����{����F{U*#��0U�)��up�*M�@�Z�F��!3>�0-+��:j�0����ƙc�z������+�n���ueRq�}�
=yt� ��j���7#�B��I��(�J�;
'�٣I��N	E��:3U�x���<>ʼ�#�S��C�c�R2�Kp}��Z��b��E㴇@.�S�S�q�����M(L�e��F`��Z��8Z�㗥d@��F��M�	g�CXsl>�_���j>������is��'�(��Z����H����̙��ɪ@ã��&�-�n��H���b!�]91g�[�}����$�Y�xA����Wv(.;�:��J?n	:���ز��BEF�� ~����I%���`�m�6��w"�d�6��8�d��o�NohY����oTXgϞ��:P>�P%X������ՙ�-3!�A��3vv!}���BTqXpv�kkcc�U"����5�5����Óڍ��r���=��5�=\K����Q��ꁊ���ml^�ЯS�>��L�E��&J������Z$�mW�,�����5�������FTg�2��rg��㩽��ӮH� ��*6(.���)�u�p~���R|X�{P��KC�h�B�ڌ?Yd]N��5�Rs���1�:t�����2z��t����0.���eaJk������h���k�CP~�P���;���_im�%��&`��?�J*�_$m�+������J�k��������Ҹ��w��}�������ؐ�D��ٳy�Cq�@Ъ}A�3�C�+m��ƅҬ�HPX[�"~�F�m���e�Jf&�\��PGyee6���r��ܲ���Q��%�*�O�ٟ'�t����a}jo��L�^��nS���5�Y�-�㼭~Hv�O���[ǅ��H�o��L���jr�ϖ�n|<Iw����}�6y@p;�:;�˟��d	�>�I��V��������9bA�Ж�]�㤫l���\@˨��m�C�.��Z�����|p��eiOܤ���� 
���w�q� �y��I,���J�ge���s��@v��ٛQ����-�oE΍�J�̻�~������f����AB�3��6v�V�#
��їt�1�i�Bx7{��s�{��j��A P�	5�	��{��ך�����7��\�'�����囗;���X��"�Wm�~E_#��>I���<P��xM������@R��oM��'%ȋ�į�� M��/}IQ�m%{�ѯ"����`��t����2����d���i�q_�Β@�p�V��݃����.��b̷qtmz�> YOEb�
Z�!ӭ���J[����C����@o�I�����d�9_�l����I��G������7�82
�#�f������S��ɀ��9 3@�h��o�r03?{�|���'
��r #{�>�$ܱ�A��tT�W��U�	3'�C!VB�d�>�����w�ߚ��F.�7R�[`��l�|m�?����<{m��<�o�
���N	�Γ���~�q6���eitߦ�ƏcF=�p���7?����n�O�a���|�g��`Yj�բ1���7ۏ<����;WP�+K�������v�Z�#�UBr	(ҟ����xӍf��틓E.N��aޥD�s�1�t@��������i4i�'&�?��ڿ�vT���9Zn5pp��^&�)-�h�����[�v/X���W2�??�Os=2?��d�m��c�,s��Jp����rxYFs�CKk�,��^�..v�sΟ���S"eP�V�c�a�^ �A� ը�'�fɉ#;J��{�_�\9��-VZF>��Nc��H���&�ƳQy!�i�BB���qc��J՚u���XZ�l]�m_�wH�|�jG
��I�g���	I8��:�8����e������#x��Z�8Y�z�Q�8����l)�a��]Dq�{�x��~Lub38�U����~EV���!�8*��R4i�hk���֛_��}��9�8�b/�� X3�%�sDO��������.�j�&��]����u�ܣ��O����a�~$F�`RKdl�����sn':�"uZ�|'�̩�;��}��5�j�-��f7�
^i�������hXc���h�h&���J���t��-d�u�'�R{m#D���r8�s����%��2vG�%;B�t���r+�ۨju;�
فW���u`jF�N&��gC��T
��>�`��;��SOl�j�k�6������0����0J������H�+b�Ϡo_��c��9�U��Uo��L�Ԯ�U<S7>�o�O]K������Uà�
�Z�StN�m~;$�N���>2w5��`��2�S�;��V��kO��������&Ǻ;So�����w�Jɹ#��i5�a��}���,JQ�2����H*n�#v�),Y�&��+�>�������	v�Ǐ[�mY�"�I9|�WD���B#s��]+���>j��#��f}R8@T�W?�,,H%�#z��N���_~/�]��z���.��\��D�G�a:�g�tp\��	UU��%2�O�+�]�LJ'��t����M+�W��tU��Z�� ���4��'��
.9,�fcXS)������Υ�G�+��hKQڞ�GU���������_鹧ߏb���4A�t��5J=+��T�hO�ɼ�_�)�����U�;#�ú��E��'�A����q3=����{�0#L}�a�Ѻ�X�Pp��$]�j�y@{���ll��M(�&s�]Q��޼"_4�=�1Ax�`�im��6<�+Hnv���,�G��2�[?���~���Jo� �i�twU�F�]�_I�A�KջY8��W��NU�5M�<���Z���|f��43�7���<�b�~F����&�-LѪ~N��>8�s���X����K_JxIߨ͸��'�&g���퐑#;vy�����.�J�Ne��#glW�{yWww��b��v���`�{В�����eS�m)h�v���r�{�b�΋r˩�d�a��������N��zf�rW<N�{����k)�J���������n�^�t ����ś;�E���+S�N}�c}������WL�ο�y���:EqmH�=�	�(���iv��A��ۉ������\ҎC�(�ra�N�� ����;����?/�9�qb���pW�Q��ж��3=9��6�\����^̳��(���ƣ���|�;���
���=J]�W;��~B��_�����S������u��Q���f�y}��hy~u��m�vQ�ڱ�=<L��C���Z��	���䉄�h�p+�k�O@�t��|�J%�0�jC�h-f�����B3������'�1y�e��/:JXfe��Iڥ�b�i�;�l��&jT��D|�S����ou�z�/����3V�n��@`�Wwk���:"�j�3M��5�^�j��ٙ��ێ�A/�#�l�ޑD`��*aJ;���7q�9�T�n�a�ݙ������6��)��d���2��v�d��iG��S�;�H4�ov~T�KV�禝�G�����;Ny4r��:��eW�!\?,\�VQ��<q�
L.3im��[�����G9ĥ��\���Ҡ�ɡ%	�I�%�Rt�@���$4Q���ᰮ�������h�0���xs��p"14/ ��(8}2���/�R�����C� ��t�S��X==�(��ld����ʺ�6�Z�A�s�_J��I]�Jz�(K����;�����
�S��'Q9��0ԓ2E{�z����/��㦜<��	Ykw<C��f�ײ��%A�q;�J.�g1�I��>��rQ肸�r� 4��,;j�ś=f�3꣊��1���tϦ#S�.ˍ�P��DC���e��<a°��d~����1�Ҽ��]	+b��Yut�U�cB�V�O�v�/n�{e��<{[P��������N}t��U���b��/%c��x�A�ÐddL}��pF�L[#6&�e8��5��a�9�5��T;�/X���.>rs�j��Z���Sk%�%���p�Þ�{�s��#�u�Jww��2��?�	�q�d�ƺϕ�������>���U�ب_,�m���6+�P-�v�'Hr������&h��5�%��ٺq�1:@�p_P��Z�D{l��� �VK�{~Z]�=�.hZ�U-�29����Zp;:�۶�]�>ԙ��8�`h�����Wj^96�9����#uB�E��,Ѭrf�FH�3r���5=�� 2֚�N��e�f�����(�i��pֵ�Z��{/P%���K�v�����W7YmY�6����c3s�<��׿�.:�+�>�u��l$�W�i�Mz�1U�E�є#���gd�Jj�^hUo���Ml�W�<�P�����C���Q�8��ķ��tbr,uU����D>ډg��2$p�Z���Ƣ�� ���sV)8:�����GN��E��:,���0ܺ3�L������C��W��@>���6zrX����*���t���Gk�U`���c�W��X�"�qku9y[&U�]���1�7���A%JY���F��=u����у�g�YV졣`�c��Ȅ}��t4�Z��r >��A��bz�D��
N�`�� ����F�cjq��J,��U�e���u��n���5������^*	�������8Qch�����8���y���~Ƚ�+��ߪ���<��2м�L(
�z�H�S���<&A\���^ܒ'"�e���rx����˯�q���S������0}�46��|��r	�mP8�gc�^㮘nT�DV�+ɕ/Jh:�N�I�9(��{�H������,n0�<�Qv�Sv���^�_�� ��=�ɉ�B��U*ģz�@a��`?����o�82��_���wX�g�I�E~Ɉ@v�A6
�+ lD�_�p�]Y�VY��"��jb^���tKk͝�\1��"t�3^�Ɯ}�����-�yA��}/k��U�
�jy���'zb�z��}Q���p��{�ޮ��a���yi��$�O�mY�%}�@�Bz�PQ��������
��Z�|��)|��t�����GAj�Y�䏰]�W�S�B���l9V~�O�&�w_��k ��Q	/�uc+L^�|m�ž-ܚ��@�����뤖�urs��;l�!w�b.�	��?C��e����1֩h���k�hG7ӂ7��^�g�Ld�=͗k�#l���8c�(��
C�m7�@v��&ʀ����ڻU��n 
$������kn�a�DOH��J��޳1��"�U��L��j�s���m����Y,��Ve|g �>,�bN�K�8�K�G?�x���q5���r��-+&��J�=�-�v)ﯨ��m����[�z҈�JأlP���,��j��X�"vKZ����6�t����V�����V�C^�X�}`�����Dll�ܤ�X��2Dv����02|!ۑ+B�Gv��r���\��v��u�v��S9�K��oS�)g޽|��o?S7�ܔ� �[�5�ؐ� 2�lm���#ųGz͊"�`����[@QZg���q��3�"��C�
(�K��/y{a+v����XGܞ ������s�6-��1�/�̴��#<��6�l��*}������`�?������~���q�Hz?��0�m�˸'��Y�I�'u����ܑ�{Q�X���n�<h�d��6������Q}	*����wgC��4NP��9s��S�n΄`�9 v�Oa'��������\:�������U7q���-O��^+� �^�U��1hg��)}��9��~��=6��'T�/��~�-�(�RX���m{?r��\e���콻e����ޙh�Lg����j����vkc�=���g�5֊�*`ĕΛ�)��8WL������r���_r>��n����)ޫ	1��w;?�����;ͳ���H�R��ކz�"Q��Ѿ��C�,d_sC�D�+0O}O��U:�<�]���u?�ȝzXEۦx��K�x3��������!?ii˨�<�	��=�F;�����2.���T�c�$�JoH|T�sT�*��=ڗlx�ͬ�H�u5[���S�kӬ��>�Ud������ّf�q a3T�U0�:�Qa��-AL0���O�	���u�<��98�UȎR�a/�ۇ���ȷJ,���3U:d���RyE �� V�%�Z���]�y�Y�w�JtP�6�̊�D8�=�>��L�s�$�Q߂*F&�v�1��k�0-�X�x�7r$���+g"��F��R��������7_��Lq9IO/�?��Uɾ�=X��ZȒX�oZ��l���U��1����&]Gs�&�4� �GOI�/oAHE�Z��U��E�.����a��UU��9 Bx�,oi���b�X���aB���K(����9�óR���Z�uX�q��,-�C�e���o�R�M�sT��W�W��al����`G1/�x�@��� �3��7�S�(0=��[So,N~p�Ʊ$���Uu�au���^�# �c��r#� ���g���z|b	3���j���J:(0�R	7�,Y����gu7��Cg@��CE�K=6%�����V�޸2���S�q\>r�	�;���l5�UspZ��Ϫ�ᴤ�?�i��B��h�m"����!�Қ����	���ڍ���H�o�3E�����k ��y%�_��P�@lV�@e��]/��#�pX��rQ}���	��0t.n��!H/�k�$�}��)�1G��sD���9�C'j��B ��g�C؆���[�	*^N��?��Mw`K�U)P��A)( 1y����0Snk�{{��#�"�7,�%��}Pŭ~�#hm�ޞt�f%h�,�/������c<>suIC}����%�����A�4��>�c���e�+C��<7��/��)���aH�{A#G�%)Z���?�q1�U��G�Ǡt�*��ꘕT����댏��lT� ���<'�a��K�*�U���� ����"[�P���`�٥+iA����g��zť���G��%9�e��T�N�e=@9�]01�?��N�)����9�$8����"��-k�����������)?5�}�li����D���7M@�������ω��\g�-��+���V��.aH����N�Ɉ'a����R�m�����Ge-b)�̔�jM-�ǹ~+�"_�ja��C �;=��-���a�g�l��^����S��*�dJ�=z�H�����X�b��^��+�N���F��'�p���=Ʃ�&�%�b���͹���-E��]<��5�ҙ��>I��ӯZu���M�^6~6�2i��%�p��B�$p����Se�|�	��4�������� �T�;�H�ة~����W���U
�z3�P��#���IB	�7��
5ֶ�Vmv�Toa���c�#��55ϖ;7��v� f�'��9!�Fb�G]�@�)��d�3;�֡���e�N$	5=��m�Wܝ3S����65��44y9Ǜ4m�9f�=b#W�&��[�DUo
c�7�+SP�h��k[���y�>�H�΄��K�Y-
���n[�?���e -�-�^I�Gҷ�i�ѦǣPq�u�}r��=��D����n�?�uKW�8ӻ�ɚ����� �֠���6���J"P���Ƌ�M�-Q���W��9crΧi� =�:��=���� �('�_��C7�� ���@'���E�ͱ n��h�{p�/�r=��ΏO�x��; �] �v��u�8U!��kՎ�l8a$1���L~A�C��q=6�~F�z����;��b��񦣮��Фw �Uֲ��q#o�Z�ڿ�  	�죊m�vP	7���)6S���sG�V�����T��=�WV� ������1D�;�h�>���Y@�%��S B�>/,�HE��!�{w}uGΠ�A1�L�%��P;���E�4vTB���g�-1��/ø���%�gQ���&c&�M�}6�5/���|tF�O���M@�p�T�0��#�=�&�(�W菔�r�KOL���23b�!l�%���k!����pkk�]�f�#�]������x�v��A<^?%�o#����D�j������U81g�>�Һ��ӧ�����Kz���Y ��zڲɭ�9�$'�u�ՌU/Ů�{�� BTug�A�cEI���x�"����Ȩ��p�����U���0�|��̱��N��y�����nІ��X`'����^`츷�P�I���v�������(�?��܌Ֆ���zl�>֫�t�1۴.l@���t����Ð�/��f�ӆ�u�����8׎W}�>z����|�n��7�osR�+w��u�}���k���n�BZ��qmp�*!�H[���еfb<�<������1��s�]�{i�K>��EG��G��;s�5Osy ��k)��q|�񹀢 ]�P���0��Y��G}ڐc?@������H��H����� ��|�z�m2m`�]w����
���Nl�Cm>����7��,���/.,��Q�it��3��Ν���b~���U��pk�5��D-3O�ak_O�-�gQ ��$,��a�/f M����� NV8���GPIwTMʡ��Z_U��.7���R�1 Y]�[e�Ic�1�04��5}����K�:��Le�gl%�}��[<�i����?\��? �R�Պ�j�{B���@g7�y֯������/�˫�)�;t�Bވ���l�zCG�[T �R��m��7�`X�%'���B虫��;�)�����>��K��f7v��Z��ǘp��y����������j������7�����e�%�^e�	ꣿ�}^UR��� ��ky�<�_	��i5e�H��ȗ9密���S2 ����qmq�˹lPx�L�顊 �._hlx7���Ўn]�2+v��[,�Kj۾�������>u��A Q�_|���NFp�V|�t�E����+�_®�� dC��8��� ����ƍ�u-<Ѩ�y��qyme�ǉй�?��no:	����8�!�u=��Е�&5{H,`��c������O���j��T�=<�H��Irlٓ	�#����I��FS�%�aP��5��4솩q�:��B�7���D�L�_X �xT�S�Wz�o���Hۜ�$��~�#�Cn�*�Y���`ϯѠSfs-�2.���"L��E������d!�C�v�fs�t�Y1�e�v���G��T��J�'�d����+�;P�ML�>�ո8��q�t)�ؙ�X'H����F�5ޣ��ӭ�� :�,y��u�@���x�@�!O�y�� �f�Ʀ⌕0�{�#[����6XA
q���yg�>o�CO����x�`������
�?�|�"�Qv���-n 6�9��_9�+�2��V͈� ,&%L<f,��Ɩ���#�&\;ʅ6��*��	ӟS�O,��1���V����L{Be�����7������E@lx�a%��>V#+�G�ih[�)���g����
���7�3V���ҟf���}�L�ͭ
s"���mM�D���@��K���s/�a�|�9�����I����J0޼e���w�r��p�?��h�u��Tfp_é��+��>4v��_��]�6�q,�6˲/��s��##G��ja�E�5_���_�,�%5���~����Ā� �Ta��\8�i#�n���&�a�@�}��^qN�8��K-!���+�����i��fwD�A�*O�4>a>x�f!s�Q���9P"B�`��޿e�-a����$�i:���=-J���ڡÐ�7_M���D�6&Ѕz��(L��7�Պ�@F�u�\M=���ގz��(GH��M�D����uϽx�ޤ�*r�)�ԇa�S�Mf~F�������+SyqQ��)Yh�5Өw�6�����bS;���R�b�8N!0���t}��+�:H�;���n�V�II�=%gwٍ�qߺ��xI"�F����s�O�E�Mp1mj�*��^�O��l���q[ Ȅ�Y-�pT�+/\C5R4��2YV��7��*Ӵ����ޜK�&$%k'�l��Y��{_��[}��\܌_�* ������7ƤL��`��@�{z:��@0�߷��R����b��Dך�՝�O�h~���,qmZ����譩�)�r�֦A�a��9(�@ͣ�Wl!��y��s< �#e[�N_fLP��Ֆ�Y-�wb�uE��i���O�kH"�z�S��|�<��@��f�)�w�a�-�A@�u�0��t�sC&�6�+���l6��g��%��쒌�,
��>(�!����SS!��q���YtSq2p?���z�_�G�+�^O}hП�|#eЙ��؃*�M>��JB��S>�}�_6n^�˨�|Gߝe<�7� ���Ạ[��'�r��C�f�J�i¬c� ��,z�ƐY%���X�3�?�ޤ@ߞ.�z$P1%�?��	��bH���E93�P_ a����v#����H|��1'�j���RJ'4Ԙ=W�r5�u�
6��.�K���K���Sl�y�c>���5���{�>�Uy�5�Z�x������܈�OjGz�0���G}����*i�Ɲ^t�� ��L�og���+~P��h�>{���m״{'�����L�œ;�V��������Oj���A����jW�D�[��\s����,|� �����iw��V�`D���z�Y��2Ґ�6�aa3��6��Fǅ\W���zTt-�t�`�\f��0�J����{DY�p�)��|�H��{2�,5���*�6��\�m���nCe慨�0������!�]��h�S�d*i����8�O��T�]�>,̨-l�͊O�z6�����++��;�N�V�-%q��'���|�:��b߿5�14��'݈+�t�I��#m�u'�Z6��vã�	���,�ukE�N�d&�����Mq�A;�*�i�|T�2r��ϝ�5�h�����m<?�T-�Ƀ��.�N1�"�S�C>���h��L�Xǲ����(��b$�z�s �U�y,�1�7>C���w�R���Љq�u'B/�,~��ɌC���`����YF�����<�
������m��Of��͙wY&�i,�.RW�0EC3!����_��sZR�
�j .� �z�L�{ڟ�1����_X��öh�\�L�a4���,#�*ؽ�>{K�G�Dy{�rj���Y	 `/�pA�������aP>u�ʞ���_�:���0��ֿ�&}Ҵ]#'mk�92��/��ND�isg��b��\'�$�y��w�-͉�M�u��	��r���Wi�5>�~l�}������ =�����=�?M�AB���.�hq(�n7Ɂ�l�Lnم����l�	��%$g&d�@>B�����̛�C�����#��ߗkM3��c�>f�	s�5�<o�Z�oi�����:Ǯ#������.C�Cέ2��@������u�+���*��f:uȕ�J�35#R�"3f���]�{� �o$��N;��Ƶsȃ.�+_̿aDB�X�%���Tx�݌C_���2����|[�X�����K5�NX��x�M���V�W%������{�_e}z	���JJ�o��P���S�XȔ� Lru*=��f�����E��\��<�.BPAOd6ĩ>ͫUGS9����m�윟�X�[(�"�Wf�F~K�p'1Į�����c�M$�����M���+&má-nB%���c�_BGx��m���xk�8����A�$���{���e����J�����lw�/8��w*Vn�{A��'��o�M���T"~R�:%u�Q�M�V�+SM:��<sR,s�w����p;�+2+e��3藏���@�-� '�9de]�C2���J^Ss��� PM<Tp�U-50};(���霒+wR4��G:� �lbd���Ξ�}p��������ʤ1�h�Z���EAR�>��n�=�C�����@0�� _ă�'�����Pԃ�M��_�6�
�olU�ݏlN�3"�$Q��YW�@�����&����2~Q4��!L��QO��(�c�ȧk&�c�r8-��c>3�%u��>�X6+�8����%��D[��W�E��pR�"Eb��2�)�@�MG�wˊ��6C�4�7C�� �����u�)X���(� �l��C�����dY���zR��r9(��(ě͊�v�w�Ǧ=�	E�'�yC/�� (��+(�-F|B����F�-����j$�|j��y
U�[0����T��PZ�H�P>z�q�t�T�:�m��q6'�bˑ�o/>jT�P��3mT�P�W��_YLS��m-�}�-1J:߁�}͝M��A�.�x���^d��z�ⓝ�f5�H��Wyo���.._˥
2Ɂgr��Hp�e���4���~�~"��7ϗ1���$���6�H@��SD��3��{�I�Y�R�^� Y����'�@W��"&vڅ}�u�`�P��l�%�=1A�#�_���+J���;7Q�]�ꉤnV������Y��E魊h�.�*��*�1���xmg�ك�w�a)n����u�Jr�+����k:TIOm�-"����x�qs���x��|�B��퀊�J���JA���a���r�>/h�b�ӕLd�HPQʅ�Y�^!E.��lc׎椴X��D�,dG(y��s�A	�PSU��o&A5�.c����|��T�MZ��� ���@�|�v̎�ޞ�5c�ʙ����?U��nc�$Lʒj,��(�z�N+'�t�+n����H,�<��A��#Z^�}�YG	O��]٤U,bpoN��D$�6�X��**ߑQk1��֚o�\\��p�n���+��.k�h�ݺ���Jmʷ�gֿ�Eɧ�����I�=�� @�C	�����q��<���87\���.��6�iP�=�	%��Uk��Z��^��=��*�c�H����1g��nZ��b�ܞ��T�֔%���3�h���<��	�44ΐ��J���wD=��/��U�~���FjqF���б恲��=�h��=��'��Dw���g�O�E�K�u��V�]�*�:��UUq!��~P���Ae���fH?V��.�R�o�k���nPO4e��F��3��Ҍ��²��/��iy���U�������8�;���-�#́ܵ�g�b�cE�ɦu�����A�
H�=@bS~�_Þ��P�w��;|kS��n|L�%TZ�M,s5]4��Dg�n_�d	cG�i{�Dﺭ�śv�K+1l-�H���&�86'�'���l�U�w�>(5W�2�:팷�19�h����#��A�S���~��NxR������+����D�x�V�K�%�NnǶ1��&��a�ea{b��!L�|�G��יp���V�v�ϵYo<z��~��e`��Y3��4V:��1�*�N��zـ��)[6Q�}�\dS�V�wK�~ӎ�x2�MWeA�c����M�x	1J���`��jqr�Γ���xL�xD$!4��{̧�Q�I䞆���|����F~$L��1h�z������帏�^��s����ٹ��޾��Cњ}�1/��*���Z��� #���5z�����5cw��ʴ;��4ua�5ջO�Ƅ���L%�I��bvT���$�v�]����^-���.�AfY����g�Y�4���=�7'%�L�E���ZDD�M6�R�*�2� 5���$Oa��a������ʫM�F���SDC}"����B�݁��ƞ�����s�<��~���8�7;;���W��_'�F/�З�F};C�L*��DB��_r������9���c1o�4-���
n'kk{�ˈ�փYN�Y�"��f�?B5os7�w�z�2��9��Y5 �4���B�<�� ��K���MZ�*)��<��D�|�<r�]$<hR��w�jړ�\��t�T"�ʛW�y˧�:��/��W@	��{��PLa�������F��6��1۔���J/+~/e%;�������j��1����A��0�Kƅۘ�k�W�&4Ǉ�ǳ�k�v��]b���@
R_��a�=Wfq`T�a3�����ڣ�* ��]O���������>����M�Z{�N8�"=e.��}"y�����U7��i�N����l�.�C�Y׽����j�����vQ��#/���:<���(P5Ӊ>�u�|��C�ﶪ����hi>�	�^�\�� ����Y�}��9�Z1f�_��-�h�a^�^q�%�,� ����٭���ۯQ�13�86W�E7�����@�#(�1�B�*�L�o��p�)�]��4���Xt\��������,�0�p8�C]>v'_��]������	�*9�ɛ'H��&������rݐ���Oi1�8ݗ]��#Z7��7Q�]��_����*�=Һ��.�2�^�=7w�@6˗K�s�ZF_�2x�֓P��c�Ly��ٷ1��{���S���a`����oh�+#������Xޒ<��)f�����[�`-�q���*�j*�1<C�jFNU` ��e�ݔ�C%J������̎Kz�������ߤ>o0FE=�Ѕ�M̓=��������k�S�@�ny
�F�(� Y.=/�{���o�i`�
�q�$�
+�%w���K��V�#@�Чګ���2o�F��{��M��c���'��O��*�=]$ʭ�wd�i�F6]����[�eWo�f��p�䤮�~!��O�|=��$k�U˗�^˝6��TP���w$F�v\����`z��B��Qߞ��Z���L�3]U�i@��ϗB|��N46�z��x7R�>��k_޶�r`������4�1�G����)���Iqu�N3����)Q�	���g�)�|�tSO��۷�_K&V�3�I�������U͡��XQC�
���~��S�z���q(��_�
�g�5����5��O|���R�!�ĕ��!���]���d`��ӫ�(����B˖�����qÄ�
��L�g3���y�~*��*��=a�K�9[�Yr���gu��K�=7EO<����V��6`|���PN�J�g�"�%��OA�N��1��Ҡ7���t���!��:d�+��->T�R�ĭn���L��~׭�jY���D�6w�}���!����$Wh�1���h���VJ�W�5A*򜫑�>��w(�=ne�rw;����-���)�rC���׾���ۊ�([��0}�F�ޛ� �֢���>,���i�f[���"������Q�-
DY�ɍ��� �w�YW��~������&�$�4��Ic}N���x�u��,�ՇF��Z���Tp'�m�1�<��{:�v���6��-�����ʢd6L�G2(��b'��xl������8ϟ�W��:[���g��pn���*�P(��=i�f�n�W<����iC���|���)�nf�o˦� ���zR�s�~bc�G�m����<���@�c'����PQ����(~U�ŠCI��i����!�r]���D��A���n$fFrh��g�����=z���{�{�s�[�w�B�SQ��ϯT�;�C #����	�u�`1L���w���T��u�n��s����JH���VM�
�P��HA��>��7L��\_�6u�A�k����]��R�E��p��P�����̕Ŀ~,ps�[j���̷be�~p��^�]w��sTׁ���{ޠ��D#ؖ�[�M��U[�D�þ�oe�~<�M��c��!F��p�e��'���lTǭ��8�����9-qr!Ի�ί�`T7�\`�sw6�>dT�g��}1){��f!-��!G�d����-��	�yFj���\�����d��Φ}�OU4�aS�5�VF�dl�"���F���͎ٗ
7 �~�B���~R�_�\�q�?����!�q��������R��NZ�����nv�v��u�6��||�F�;<�_�}��J���Kum�#s�P����o��Ώ������EҖ��m��F��5�0^�Z��;?�����C�4ee���^ca)a�-(����
�>��x:j�"���:�(�$�In+���2�������?����J<�5��~�_d�c���0��m�����c˹�2*U������U,AXZ�/3j�PݵIV�V������˿��z�B�=��?R�o��'�1���x��V������R�ƈ @�l �\ 9���)�ǲ����ߧ�\!�6K�Mil�<���a�d���������_�b,t����݊�����,�qqi�AN��T�:��4RWj�e[�{-c��U#Su�l
�3�߷:���@�]L:u�����_j{|�r��{IIK��K����)�А���4A2zz	e����J|��J+(PJ���w���VΊ�3�ݾ1�*���U=ˋ����~(�S��q�}���E��*��<1Da.f����M��*9e�>}J�ҕ�ș����ޝ�����c��@����ǻd�;�j�?߿NN�*].���Ƚ�%�A�\���m��d�\�k��^�O��&�G+��ׂ������F\��+������<,ƴF�]m9mL��ϝ찺�BW]7^�R�z���L�?��=&~�^�8/-+'׸�j="X���k222ߗ/_R��s�7�d�j=X���0���
����`ؚ��1W�n���nN?!�O�dl�����:�����CV�{R�׊:&\�&͝0]���Ls_�c��ܿ�3��S~5_=;5f}��Q�`����f�\�e��X�v��~���̌a,܅�]�"A���h���Ԕ\Z:��ܥ�h�S��&:۸��\{�noc�7�zC�����e�b_׏����]�#�<�L��]~XO=�a^�W��,�:��>Y	L�՘k�O�����U]j��
V#����n멌$���F�9:�|@���f��`0��������)�C���������~��e���_pkO ���,Q�>��FY>�>e������PI�h�v�u��2o�i����aVG]�a;.�CH��C�cݪ�w������*"	A@5L7�p����b�b˨��F-t3M�f�!�* ��^�	gh���pQ(��&�E5w?�����߯��K<^�4��!0�y�nO@��������x�y��yP�,�>�:�H���L
��Zia�Q��EX]���U]Jѭ�����?��ttt6v�kk��/��Od�ſt�W�B���մIϱ쵱�uO��]5��6¥�������*m�P�g�Դ>��ܧ����r���l�
�J_D��.$�ē]�=�f}W�>��연3o�QTTRRRv��2;�o�),���j��!I�����*��K���lT�^E�Ѻ䫠8�jU��um�|�,�\o��6��O�G�D �e�N旦���o���3=��(*���v�µL�j�x�_�Eʈ�en\"��G��q�������;�T��ml��zǫ׆is�B&��w��s��\f��O6K�����a�i��5UYM�(��sZa/�no�K��<�L��8Jb��l����sE�4��r�Z��#?�,�������4�5z�mvҷD�|�v��S��2���hwӊ~_����LKL��[�3�.����+]���55��>ZL[���}��R�m�5L=�ȳӎ�4�^*D�~Jl�yP`2L���W�����S����D��'3��6Q�2��\��7e��|4����J:#��E�|�^�3��6�����M"�0��6\fc���+V�YZ��c-6�V
n$Y�m����ũ�����2�����)\��l�<�1p��Xu���y*akE a'�;��l�*g�	�8I����o�.�`2�`</g:u^��M���є��+P�C+I�����7��L�:[��A\�;�%u�p3a��O)-�G�5���ا��C�0�V�$������ɏ�l�'�+� �4
�QD�m.���	A�l��e���K�ʺ���2�&��,���`��5l[q���a�\�������/#T�nb��f���kl�&Uܘ����,�f��;""gB_D޽������r�H�F��g���GH��Uk<�!��b����9�4v��-deq�e~sJ�RΚ/+��/�f��?|Χ	�����9-�^|u��5=#���Mu�\p�g���'Z+Q���R�L�?a1>�J�~/�g�^y���?"X�ҝ�.��G7,�5�d��w@.�`�E��-C��)�io�ʜ6"I⇊�b��<�Fr���b:j�O@��m����J%���y||������3�L�F��^�|���i��&����=�Ϳ���J\GM�S�0+g��V?pQ�ig�_���h���;��q80x�h�oX�|kk�q�����Enddd����fz��=��FicxZ����d�>ܲ�kέe�lC�b����� ��'��)���`�	�")����=>N9x�;z�z�]������W�T� �_�i�����������.��yg��^ݟ�'��͉k6 ��C���.,�����J�;7��闓�S��I�,�Nwc�4�4!�>m�Ld�u[�K�J�F,O]�$�
I��3�fQ#W�t���h��N�Rf�e��$I�)�����n|����:�����j�Ը:
g��8ب*p�J�a|+Ek� 34��t����6�ׯ�?]�[=%00���(�_0�����,;/ݳN~�r�H�n+���PI��1�}l��tԇ�������{
��������`��d���ה�����/�`�" _�2666�y��t��N�QBoE������W�Zw
�:�P�?�N*����0�T��Mc�uF:��Jί|h_�9�C����,�D���@�Sҁf?�Ƅ��F�7�Ya>ow�ͼ���y"ui�nt�oal쟭H��~G.���v~��h�����C�N��/	M��7ސy�п�eY�3=&������|�ĳJ,~�"�P�sz�ڇk��6���J��c�N�����:
}VM9���4�r*H�'y��}��_1��b��M�&�Y����~˰��"n}-M��3��T(�3���6���H�٢5�@�C�+*��8o�u���3ɯ>-/�Fi�_^^^t�o�GY�������z�h�^31q�,W�l�e�'b�g٪)�Y�%$Ҕܦ�����+*(¥�_�Nw�Ǿ~���jVp�+�Ib�8}���*�QR�����GE�ŏ��� ���dK4����o�7����3E��WUQ����\ooo�3���{G�����\/v5:&�|Y�]�^*Y���|u����åɠ�ak�����h����������M33��|�N�m�N7=�0�FOfl닳�V}D|��\�%+pqrz�kV�!1��n��=1A�B����¥�܁�~���$Y3;]��Y��C���As�����6�VXb㗜�����ގ��
����X����E����W�u�jY�� ",,,�ڲ������klۄr�%%�k��O�>yF;"@~���_=�� ����q�%\:��_*��o��K��/���ƴ�߿��=�ؙ�z����o�(e�::r��ӟ����)���)))t�Ԉ��Ŕ�\�����35.�>�� �~��t,�u4�ecckL��L,��>ܫE��ױ�H>U5���"� ���[�H���#�]S�@z9���9�p�bM���M�{N���S�\�9������6��ϕ���xs;;�۬����?�����-���-�U���]�g�-�H�#^����>M��C�G3�;�B��៕��E~�ڧl��D�?�����b%�5����<v�k<��5����&&&~��ʞ��vҖr�|�ׯ ӣ4����)��:\�>������ً�9	�~��C��/&&:�}kkk�����ƺ:1�o���OY��7n8�ϗ��~��̈+1v�p��&��S�K���p1��j255��@b��F?�"����#���]> �x��'�Addd8yyo�r��CFԻ���}����Qd�K�����;E���8�H��ޑё���;&�(�s�hA*���я��Ԕ��B�ٱ\[VV6��]��M�%I���+S���9ʁ|���C*aa����z�랞�� r�1:L}�=ql�����v����576h�5\z�9�E*�'
���[���ja`�����gv7�o	A�p9�X���<�h�*m�Y�0�׃�A�h��'g�M`RRd}���"��{;�%Ξ���^��j������JS"������A��bG����RQ!M��6p�cY�i9��^jlL��͛�R!E/� ��2�x��U�F���N��'�[�e����\\��[�{:.1��9Lս���Th�i��XAy�����`u$%�M�7(�[qqq?��>G�m��*pH���'�>U�Rʒ����i�sO!���63��A�ӝ:QB���U�V&,BFA�~mm�Ŵ0���h	�D�ѐ˸�(���M���W�pk�w@����NT��7~��#pp��o��3���	�gY��>zm��	�@���+Y��sq
	Q �;�m.}����n<���o��5��� s4B�>���HB�	��c��Y�VZzp
�O	���a��S_�63A]�q�B��`# �l_�r��C�o�����z�JK��ㅑɕ��Kf⅄׮A�,V�S�2ګ&���[W��t*����)}`8�{�" �����F�aF�˗/<[g�o6���!��	�6z�KN��$�Ȳ�&���Q�D�1g������� $ i���d���襢��ρd��$����N�kjZ��	>��~��G�bv�0�lP���]���0鴲�7� �*�\���oje�qg8���"\XS�'�F����kf�<�i@����._�,@Np0��`�w��U��g+m=5Fȝw+E9:��d�tw���4G���n�z��W�D;�����v<�]z��)�a ��eqL�Es��+�djY���� �Q��>a_lQς�ר���r@s���@�L���B�/u�f��)���M���EIE�"��ׁ+�|�>����%jv��0jp�_c�QUtl�(���ɍ�>�-��(R����j�����$\���A�433�p�kY�)޹Aҋ>#7.X���J����^BT��׃hd���\���ƩF��å �%��X���0���Մ�T�ٶj��'�;����s�oN�H^�oוl0��h8f�@�=::����m����ίi2jj����I���砓��Q�},&H��*��Tȷ�J�SCh��oI����] R�ӽ�u��WA�.G������9�f3v%��{Q��q�	b|�����>��n�K~-�U�r6H�)�L<�� �
���w�@�iθ�y���[�g�^�'>���`��[+(�{੕v-��@&9���� �·J��bnc��5�.7�~$���4��sb'GO�*k� ��_~����5BAP�7q�s�'��#��{�>������mB���*�4.*���Ċ�_��7[
H�<v��k�_��B>~������`;$�M����u��R���UmYY���`����Q@ �;�3Ȕ1W$�����N�����޴&���~�@�99��; ��uƿ����E|��i�<���׿����z�Z0��� �Č�t����͙
���^t
?��p|�X>i��x��ѕ��0(�l���i�TV|�5���c��>C�]��dR!<�
�A꺺�gI��v�4;tk>"YFs�҂�~���wڹ�����1�a<�D�	��\�̪*����_K1㕃e��}It������r�>��w:4�����Q�K� ��]�FVnW`Yly���f����;��\�?�J������.��7���OЀ?�~�O����G��N*Y٢T֠���W��B��P�[���OБz�����M�� Xp{ХN[�꪿��k�x�Ĝ<<7+]0�?��s57�ΟP�y����*i���GS���D<��:`%	��QRZ�$�qL��!�p��;���u���]�(d�F����:g��ěPut�!2�&��3�n@�N�=�{��.�������l�b�I&)���m�sr���P8�$ZYY$����!O
�H�(@y M��g�V��F%�G�a��,;I#�C�bN7SeDó�vbp�U/������I��w��V��"Em-��K� �G����L�ݴ��b�?������\Q<�7��-���m]8.	�⯧�|�p��K{_����\Z\���R��V�Ύ+�G�j�cS	�����)8�<��9��6{6ZB�+"_F���m[��ek�n+e����'�����һ�J��X�c�j�� b�Eƿ��V�� ��0�}q@�$ص)G��3pu��ǧx�!q���A^>)j���pv����O���l3֣�� �JtE�4�y!7ܹH�~-��?�B��yu@LN�!yz�Z��;�cV�����:F���P�t�u�IO�r�{�����B��g٪�^����*}�Vc.�_S�-󎄢+___��!(~�Z���;�94S��'>�K��O@(�C�����'�/@N6ttȾ�`]T$>>:��j� �j
@��KU���=��p����`�g�p,h]6H�t6����6:@W���$~����^\�8���+\X\���S؊F
a����T��]��4Ֆ��gA��LZ����ozz��8zcdX)��/ � `[�E���P�qP]�իW���ssr����M���~�4m6a�4���Q�~i'�t�uB �Y z���]� l�Yk�X�ѣ��s5�����ٙf����3`v#�?8�j�z{{����.��
e�  @�y�f�=�3��N�e���A �y���y(��.���?o���0d����M󽏏�6:� ��nYL�W ���`� ���XX�0��pV(�>;f��"�pI��{�w�#(����t������HB�Q�e����?H������p����l@�qm�0���<y23V�BN�T3�	� f��H�7��р��0]9"I��(�Z���������\iU�A�3S�| 6��!�%�0Hb@$LVʔ(����xzoYm��B��A����# ������v�*{��#�Ė���+�K��JV?�<T��4p��]'��!d������ jM	�3 �E�>��#�Q�5?=���}���uǳ3_$�1�Ùå9��9����o8���rx��$-��05�mK#�0"2��As�݊�5��e �L�q�~= v�N�=����e*}IYY� #=0W vH	�����oZ�Z��	�g�UB�-WX� 2s++8�T4H�oD���O\�1�vzR� �1�/������-.)�P��Tw�"6P�\X�}֕3�+כ)))������h`~'~�شB�"�j<HuE�>	���5����@|�m���������/��_�����D���x�� 9Ъ�??�=e�zNNNh�Pu���/㢑}8�&?d�)8FN�qW����x�"��&?<<<F}���LI�G����� �Ƚ	N�X{��1
�|#�T�=AN.u���q8���(e���� �I����ߎ��
���'�Gh��l4�8�;u����Up�'�H��9D��?��@���O��!�����;�2��P���A��Q>��5�s]*R!�����@ �{�2,B6���V������d ] ?��}>���j�nR�9��ܓ4��|�'Tq7�UB2�m!���v�D5b���^���w�lq�����~U7�G1E����jMa��S��wf��JU�k�M����
T�:Ju��V�e.���?g�\<�D��E���,RhXNL��H�@5��������dX��o�?�|>;��oƚe���>Ig�Y-����$%L����oG�kC�4����h�o)�]J�kw�.�P������Z�D��BK��"�IgC�bN���Q5�4R�(,�֊z-�b޹x�W;x-(�XĘN֩,FV��=�#�`h�^n���1׺K���6�m�=�[�LpU��ƷE����o [_���%#��}Z����x&��֯O[����]�/f���tI�Gc�3q��ލ�؉��M��Q;ݤ�|5������~|�cG�:�k+zǯ��5ۗ;-j�R��-��i�_��NArzeu��s0��{hҪ}~��s�����#�eI/���L����+�)W{C�x�D�&����VOG��z�h�����	m��ե �%b�����z��$�3�u�1��0�DC�}@-z{0��m�[��O�تt��>��������]�x�P=�����Q�i �z7rT���9�7�%��w���R����yRk������u1����~��T�x�`����� 1��ÆB HVaI;��c�e�붱1�t(��Ӧ���������\���%/�7��[�������b����=�[Y^~���P�8��QBO���ڃn��XĊ�~.��tŸ+�oY����6s�moo��=��=v��8 ��� d���\U饔�[��������$6�ik�gf/�v���
�Z����������˱\{s�6ۅ6d	-`�gf�������+Ǔ�u�\�O�F5�v]�ܪ�r@��������y��t"Da�\��=]j�p�@��5nr�*l��@bt�p�(��?��C=�ֽ���{[�E����N���G����j�)S�>�^��K&�d�W�"Iff]�_��`kЗ�+�_4�f(e7ez�9:کm���T�������{�e!%����}s �o���\���Sz���B�f&=�bf�kw�@��?vЪ���%��M��A�Ӏ����*���At�q����j;�g��E=o����E۟F��kׂ]��h����An(I�����@����o؇����%�klH;;�&�Fڣ����tnlH@|��2UΒD"�z��C;����'ڟ�%B�vk��r�����q_֬�Ȏ� U�h_�ՌY6�n���@n��hv��7��M�p/���H͐*������$�0�C{�JM�j�M�����_��m�+�Θ6K�����5�ބj��HR�>ĞaՁ����5�a��h�0W#�F�v�FG)��9���`rz�U�m�&D$��s(���[�q�$f�|y�(.)�e�+l�*����c����ît�ÞKGHL��z4f�~ѻ!������srv~�#'��%dk9���j�!{�~�����u�[n�?:W��r��� o�	�n��c�'����ǈ��
w�l����|����	@�ѐ!��KU=�}����uϯ]Ci�ny#7��h$X3����hVcv搳�	RᡠjL���L���L)�ܞ���� ����8���>d�Y_����C]x>{���h�6�Z�`7�M1G�6�L�y���S	G{�h,t�)4u���!�TSS����ǂ "0�2+,��i�T�7�5���7�)�+���*�L��F����l�ˁ����6�'f�V�8�)���$4L];�e�n��-� 0>8�9���K�z!�eu�}���H����q͹�A�R��Eg�)��Uq~��7�}'S����OL,q�1.����i��qV��#��/jl��3�J8~��=͸�����J��ᗤ[[��X�u@��5�o����m���}W��H/�1�/�5�ޫ�ܴ��.q4���:T�u����,�xQ����}����d�O ޥ���.k�w$�z���<G@G�L4Z�%���� 
'�>O���%
�GYK�˚��_?Oo��1��I��V�"��Pf��~�^�ڞ�^���є�7�Y_�'�c����\j��&��җ�E��e}~̿�=��{��%���D)�������&T��C8)�P�n�<�HL��X[�=�k�K"r @߀iJl�v�mq���<Q��e����?�A
���j��s�[Y*Y˲�A"��g�IR?Ǒ�>��8��8l8�)a�i��,fx�@PtR �Low�����M��Cl���+��I������Y�!� �JZ�|E.�c�/���N�1j���va3�J|+57�2ߞc3���ز�q�%�}pv���7��j��Z|k�fM�������c+�c�;;[���RO��b�,� <[���	�L��Ų�����mD*<�p�c����+�ȑT�s�H�R� z��s��������𮂊�����B�͊-w�G[�Q���B�#~����IVSI{����͓h�A
|/[�������s�'o�&��vm�{��E��F)�7~֠[;���+�:�-���&���t4?�lk��p��`M�L��~~2�&���̖k� ��qC4�<�Ѭ�n����V��p;!�f�6���_���=k�	IIIHR�~'%�<��5F*?^����b�����ir�{d���q	ѱ�%�)�B�^f��W�`w71v0
\M�c�s� �1Ķ���-Q��0�hrrSX���'�E����qU��SF�D�+Y�_���'�b���{�h��$�jƊ����&��1;7�	�#�@�-Dc��oK&zG��
��PS� C2�����4�ʍ��D�K�VG��OCR��=F�N^��`�B-���B��������8�X+0,333 j��������S֌��?�����
O��4:n�M�Zl)!q��3��N�&�<���]�f��4iM:z�v�׏�h-]���^��z��Q�N(f'��t�h���NK�D���XS��}m��T����.�|�nm���j}*�II�1��Z=+�1��5�_/�����"��-�b��v������M��$������jX��.
���o}���m�CLc�<�V=�u`:�ںjs*0n��GO=��Gg;Zo�L(/mD��q�k�ۥo��	Ōn��(�r���ʽ����7�{��碳��?�9�ϥ�Pz�6�8��������#�:d�'���T-�)�*DU�P�̱�<GAO�f�.=콟9����s��լvwA�H���6�Xu]��6�F�J� :�(r3�rk�y�w|����I/��me��f��s����C��9���#Z�IL���I�;��r1Mj�� ����8X^�N�ޱ(Km����}��P�n)��mz�sV��w���U��y�Sa��Ϣ?׮���,9���-�/���t��S�VYe[�Ń�:g�{�cQH��R�����C�m�3�ۥe���KL&{>��(��q�픪s�;��U��n�Ţ8	�tk	6��of��{?����h-��؊���j��QMp��g@W�K����	�p�e�E�
ͽ1zz)G�v�$5�'��� ��-��d�,%��?�m�D�D^&�s�e n�iZ�˂��x���I�(��;QsD2)�Yq��ͭ���'�
�D��|�~�h[���kL.`�`��uf��}���}?k=�2�ܦ׍�'mєG2G��
s�Ǜ�R�=���<Q&=/�۹7WE���^���&
��ri�ݯ$Bq(^�����F������*���l2�[j��Iy�|	�bU|��q�E%ܢ�9IS�
k� ��$�r��<w��������8"Mm<~c�b����Xg{m�Y�����z�H�I�Q��G���f���	��³w3���iIH�xm��y���伂
�W�?(i���G^Q�d���+�}��P��>�*G�O���[\��~)J@#­�������(}$Ad���U���&W�tQ�]��G3���}�������z@TB����",���6�`��Tj�L���笄I99�.E���y6z<�8���^�q�#>��[�9"4���0'�óck��l����b)rB/%�}�L]wF7�F�9�QL=�����_p�tn:�ˬ��S��`L������]y����>����YWA�q��lS	)�u�o%YFqy��Lz5+�I��_�	��9��&7l��!V��6#��7.�b<W$�U�����M�o߿��`�<U+���/����h���H�QeV�h�[��������!�A�s)�>Z�
?��j��t�d�XzC^|��[]Ʒ��Z��3~j�lx�s�\��۝֠m���Pf�E�c���\�c�QP��`���.����K#�x�5���%� j\)�z��U����a��:��i��H9݄���g�sH����:q	�5�7���3�����{��*#�gG4`�� N�XS��
dZ�gy��Mu�U����VH�i�2��̍����"�m�dnv�����
�qp�<�D#��g聈Kb��:�	8��?=Ikilt���ȹ���6������Ԡ9�	Jm���HDy�W�R,HB���0~��r���,UAe͡O,n=���#��*wv��ԏ'{��t�b���z���3E{c8H�@��N<ჸ��=���x;nPZ���u�����J5�TI�I��p�aT6�i��¹��Y����O��֣"�{}[�}�>I ���A >�j0��2ģʢHE����bn�h��0���3Z���]�y{n`�[[�X3J���������ZK�[yp�S8��W���c�!�d���ݶSO<��*N X�Y^���i݅���
q�B݇�d9#�"�I�d��Q�u�d�j����Z�v�#�nQ�b�Ŭ�U���	��_�	��/����4������`�}��/v�,�]T�ik�nJ�#��+�ƋJ��H�>��Ӕo�Sέ���=~��O�p�H0��ll�8���u���G�W�2��&���u&k�Jh6�C��v/��������y��:j�?~�ϵ70�qw�j��_̎� s�Z�a!����c{�6��h��\�'i"^�5��˜�
�^�do��"m�1�^z�ax���a:4A���7G�O{o��|0��G"X�����X� ��+$:2-?d�[j�+4���n�Dy`��_1z�-ҺTx��c[ݔ�C�y^}��#��r��9��9��l�[���o\:�����v+�y��KE ������]LQ��Bּx ]Z�l��9�; �1E���&P��H�;`E����o�&�#�ݜ,�������c�l�W��|��}�I�e�6B{=����Hf�$��&��휘w���#�Hi{Eun���ư�^t�(��԰���KK�k�԰��C��^c�5h�ݛ^G/?�(�#洿�蔡��*��5P��`$c�[-m�۶!�y�\"�����X��>p��%h�#譞L,f�]���`���^u����������j���]�%U��!����sƔZ#��^��7UZJ�u��L4�p��T�b�]�SO�pcU�[���L!`�@����QZ����Z9*���uX2��]���o/��E�Cw��L�����>�{�:��R�@:��E�`i>GXIʆ�Ҙ��`�o��+�4:Ô�_3�5g���?u��������й��E~�s,���hN��+��8�j�7b�y\}����r�5+�%�T�O;���RA.�#�����B*l���S,�w ����X�wy+0c�#5T�C�m��ƾc���Aa伄�|�������g�º���Rp@$��������/�Dϭ2`u�3Q�a�+�<l�.�x����������=�IÈ�J]?åG믧g�}7���]+�=l��_�x�>��{zd|�����+��+��g=��F\V2q�Λ��@�6v*��+���Q����z~0�i��)잁��m=�&)��)�X�������^C�g���n|@��\OvϯG�]�r��Xh��a�D9������=��hhj'�E��^�3��pMІuRr�@�UxB�æ(�COɘ=c�A�s����"�"��k��y&��wv�6�8_+�?���ߡa�	�Ez�� q%}�&)�ӧ_���!*�(~�xh݊��47�<闁�ϟS����p����*����	ˆW���S���ёm�}0�w�\X��V�|�gM�+)6T'\�p��)���������a�O!�d����tS7� mT|~��#z0B�@|�+��<{����O>��Ͻ
7u�
�}k��#�U�n�v�/�7Of��:̕Zo��f�b�}�������P��Z�䝒�]{k4���`IA�� ��z>R���};��[B�7�aN�IA\�j~j:�(Ց�jJ�n:��v�CC�	+�Q��76�Z8��&$]Q8���z ݑ~mˤg?$��{z(�'j�o��Nmd�5>y8�B���-��"-ک�'�m�2v�����ؼGh��/�_�W�"Q0܉�=����@c�P�?�9�74=��SO��f�����]�L�ޣ����@"�V���1�J:���+?0/��8�/�[�ܧ�O{o�{5�^����O���$(���8��\2cxu������yQ��$��2��
-!�#A�^�)�S�������sǭU�4���xd����G[R�RUp��O���+/��6��;���u��|q(�MYE�GpC�qP�Q��9J�U�;<�02��J�TU��#�ǘ\�L�}�dqȿ��	�Ȋ)�V�y*)t�A>#�F#O�4��a۱5[e�[:moǽ���|){�@�w��i.fgZ�;/�^w|K*���.�:���8γ�RI�]�����w������.��{��Y_H�:��[�*�%~�(vy�=��2�u��j�e���-^!��Z��%��6���{�����u'e2�F�F���Ā� K�sݮmIk�ˊ[sa���k�p��*�6�m�t	����8؉���h����T3��mc��|�g԰u�$p7�9�n���)���S_n��ʱȅ*�����'4t��:����ò5�#K �����
�JPԴe�x�Y�����؀��r
�*Ļ>���˹�--�����5�\{�f��Q1յ�\�I��Z���}v�5����D����K�&V���+]B'����m�Q��1�B�\�;�A���_���,P�7�'�!�q�`L^��`��a�ZE��U;BNU�`��ff'���S�{�FC��{3�tWbl��Vx�Y��^����x�'-d����@���R]���5%5,�a�Q�}�la=��ۓ��w��Ze�<B	4��7��L����'�ٱ�%��퇵�|��Y�c`����uq��~:R9?܂{7�:[7�;b�{�9Ɵ�L���\1Tx
"m��v�u"'��zޫ� �.4�����z@p�s��;uA�;���
4�>����N��������׺��qs���7��BNb�n��j�sI�����?�e�xX0dL��5�ͻB"6͵�m၊M_m�jU��^��&
zж3*C���j�k�u���_N�M<{>Xf����ͱ@�*$�������ɬ�Z�X�k_�z�]�����5]y�+IUi�:D�K�=
R�'���h�O7>��+����/���sU��
����1�W�^�U�7hg���_�J,YBo�Dd������!��mX17��MuDW�.�O�S�/�����?{Cv����*�s��m��4��?���fZ"���N3�2�:G����+!����2v7�8��J���>	��%�g��B�^i�\�~��fŸqo�o����gW�ɽ��j�ωt.�-\~��V�[FyѶ��ho��N�k�[�o���I�<7V�B=��v�	G�v����_�o����S�!�_y��U��� ����S2r�b;���W�M;�_ˌLn��C&�IW��mw&Z��ϵ��4�C=�!��J�\��E���C���Mo����p>�}p����'���7��BD�:��Z�������2����{3��hܩ�GM�fX?�s�R�%]Be��߷��kr��"�Ll��GNVz��Xk��N=.�4���'�rh]�\)V#�Y��k�����\��[/�l����$�7��>]	%/�ڊ�e�jg7����N�4��\3<���]C� GM��<�ͯUe�D:��Z�����&I8��%[nUm�ƿ߫��f*H2K�{�8$SK�ߪ������?:i���^�W��b�j�e�qd%�鞵�H���~	�C׷c����M��v���x�A"[K�Z������ɽ��R��u�T�Ӟb��J��*�μf��k!a�}�M˻��S������p���vF�n��J�[�5�����>����!�VOO�D�֮���Qm��6]�����Zd�.QpJw�����$v-���F��ˎ�\r��t�7{�zZ��z^*�R|�ט2:��5��9vd�N�z�>�Sm�3תt�	W�Aٿ�7��Y�6�0F8����Vk	�����O�DH���]���7��1�������.�A������+2���*�7�P��ގO�ꜚ�h�Y�ֵS���F���<Q`sO�`n�-�I����/��V˨�?���z��?��s�X��A':�/�Zk@�U�Zߣ`YZ֝��e�7��[�U��,��JI1�{�9�Q��)�^����Sn�펍���$��/A	��L�w6	ɬ��Xx`+Z�Ǯ�ޘ��`_�͐>�q�?��^��P���S��!��C�K���&�$�薊��=���WH�4��8O-QZ�H��,��z���^c}�C;T���󊫈?ܷ�f��V���#*B)U�52�c���1�g�-��g5>�7?����{�tt�^(�;�1�%�1���鐷�Zҍ�~��H����:#H���GGu�Ũ�����E�~�MU��{`���63�Ar{���n���n�z>^��v�^���)����	<�a���ݑ�q����ž���~�L�;�Ą�`r'�hHw`�v�C��]�yiXtxi�����s4$o���V�������Ki���V�VǶ�.S�w��Z�e��.��`j��g�I0�$a�o�NV}w<\g�-my#<R���r��~̀�����j�4�w��UlS�oWL�J��&?���\`x8�g^���t��r�⤜!������j%��h�@w2(�F�J�9��MSV[/5���5Q����A���9��������[��UH��zZ��1���Ⱥ�&����DiOi�ҥ�bA��ҋ��� `�J�EiB��@��ޤFB�bH�	%����S?��x8�ν3w�73ww��u �zǱ�1D�Y�N�Us)��`�m��=v�����[n���"���&?-j��Vh��	�*�<W~�<��?\�4�@��X�W}��r*���F�S�������%LYr� �f�ȸ�3L������.��2��	1揍�������e��Q�.�����)�m���qhӾ��y��fV���*cm?�����$p���8ʩ��n�i�o(�5M#{'�0I�T���#Jo����U�������(�z^nPY�L����Du��[�a|�?�:ĳ�,��r�$=X˝�6֖�p�mT�ɟ�S$J5J�P���ޜ��ѩ��4��cL2�P���q�[�s����h�>c��r	����������#��������UW�+V��;�"�M(�7�<�1���X�|p&O�c꽼��a��������/����,�Nmۉc���R����F��	�_#'�m�Q��yѺ����;KM�����W^vtɎ�H�9���"����Џ���{A3P7�}�W�R=���H�/�c�ޏ��vp�1N�G��yW��ۚ� #�E�Հ.�kS��'<�#ɋ��L%�~��t u�)��>4[��賿&��$e��#�v��`���&1]X_�e�;ѫ� �S���.=�>�ZɳLV)���z�!��<+l���t��|)d�)]mՐ�
s����m�`�u&\�j�q��3�R}��;��ѧ#�D�#�2���j�cA&�}���i	j�14h�}{�|�Y�0d�	?,���G5Mnƒǒ�M���\3|�Q��X������ܙ�?.����MY�|; �� �o?�;E���$��ќ$�}�0$WS������'��H����e�޲2������5���q���)�ma�x����8x�E,�A�/�a�"�����V�"l��B��L�'�P��p]�U:�GI/���N�U�`���x�-'�Ӻh���GGz~�=X�a}�J���� ��аo0�O/@�*P\1=��pu����}�i�: eӺY�{;�����@��V�H��&oK�MY�9巂󬒻�O���A���骉,k��x/I^R�������i�L��m,�g�;���&��B*!�
	-ͦF���ը�x+I���	 2��-b����4�U�ᄹY8�l��&��Ĭ��?ulw�p�f�Z`-�(	��|���Sq��!+y. ��rt`$i���$��JG,'���p�1\�~��cIY�����&��G�^~5!z(������7��8�&�88؝��,p>�p���CV����ek��Ks��$�mH�m�@���!� ��:px�MBl�{�Ա)[���׶T�=�񟉝/Y'K?��� #����U�f^,�d>���+���f��V�1�����U��B�����4����)���z+|��x��crN�����"�'�������i�T��_�7��������!���W���������ݞv�5�r�Oώ&k�g�Mp��Լ��)$�-��f�d�=����{_��$t��5�̬�w�e(�k)������I#�����]w�,����.]1� }8Pn�B���#�;��
4BpM���=��C( A��A�>���� �)#Q6w�Ք��O�H��,����Z�Her�ʈM��GS��� ��&��y�8K�>�����glu]�Nc�1�י�TGk��V�DD��wPIL�%�G���p3;/IRj�cIxu�*��iu}���k@����8��B�����K	K������dZ�"]ԕF�L�>ߥP�����gc��@Ѷuha��?8O~�_W�<��,k���J
�o��������̊n��T�ɛQu�̸Ք�����6��Jd��=D����R1���~��H�����C9$-W-P�J��B�D���V�B��4_�I�Y,�e����_I�`�I�}�|K�7?3�藄0g�����KQZ��Ő�~���� ��z�E�%\-���_60S�4A\����zwf�\�wA.]�-��:Ghnڎ�36��#	�=��{�w���� Y��:O��;��sjӓ�чr�B��=đ��K��7�AU��Eoi�,��{,:�4�_��
O��.��i�s����	b��Ey��M�?),ˏ�h}�^M�v|�s�;y$G���,���-����1��c6@"�6r3���f"_p�=�n����C~3�v����?��m�_O֮jrsS.Tm���Av�j{�< ����M�^�3[�9hi���Kn�Є����#��"�L#��I�nmE��};wϻu7�v1'ϵ|B}�L�e���m����ȯRg�2,��&�Wƺ��͟����[d�A��	�9 Td�F=4����j�:��ma��߳%1����ܐ`յ���
�,���9`��pm��>�DW�I�Dо�V� X:��O�GɁ����������e*�:�&�A,Ca>f�\fKJ}�w�~%��8��\@�W��U��$�U]c���_Yۀ�N�̅X��x6eU d��*��A�T��ٟ�W��Y�\5x�Gn&j�S��p̶p�1I�O.�]y��L��]� O�z�<�X���<�|�� _�*�� �F?�y���5��F�6�LM ��=�����~�Ќb�!�_g3���n,>�D~���(�J7)�zz��q*��q�fTkV/�z��k	��q�TfY�k�j�]!>������3���;��_�("�4 ��{|�j�x\�eQF0"l�z��Q�M9oJt�����RM���F�j�\��]�Pf{q�rS�e�ͥ�:�w�\ߪ��u�Ў#*��
��iċ�:�й�k��'h*�� m3�E�~k����
��W35�v&��ՠ��tS��5xuY
��LB��s;W��~r�bsn�*��	��)�u򚒪]����Ɵ40<={��2w���D�Dи�r�a j� �b����9Bl�
B�N� ��Vz0���D�O���J�-d�-nz���z�C�/3�b}��},F�{](�m�ȍr�͠��&$=��]���1o"�C(��μ.��	c�/r�ǚg����yVY-�9�Ǝ���5]6�|.��	�]���^�LqAq_��LW�ӹ?�=�V׶�q�o[��MUE�SV(ࡩ梪ôcxwqKȒ��D!r�7��n΢�Xݛn\ǖx�b Lo� �ޒ��]^���t��������Q��T%����߂LU-q_��2�����z�<�V���R8k]�J7 ��8i����ΡN㱚Bgc�ܻq��߿��癟�x0P��p*������5rn��c���J�����5Q. @ ���f�6����3^��<�hBR��d0�Z�#���et������]���G���DA���qn�6����{�!��ަ�(��n6��q�^D��B,KꂡC���ԬQWv��`1��a��'�!�ِZÎ׿���aj�3��]���r 3�7�>xo��k�U��#���s[���D�\�	�QK���~��t�P^i����d����:a��.Y�]đ�6�h'T�����߂�#������$�I6���xs/��O��7��@W�WR�{=�@�2��lz�� !��}Z��q��Q�#V-)���D倨��!���$�sȹl){�$fw?����� ^} O��䫁���ī(ҕ�0˙��ܧq�I1�Ǵ!���2lLU�h�qI�v���v�T/�=�]V�I*�,�X m�k��'����F�tƠ˝ӣ�B�Y�8�)�^����l��Lm����U���� �ء��B�dZ`L��*�g֘�Y�BK����e�C�:�+�e2W��
��-R�&<.)Y�	��Ȫ��A���DP՟H�:�52<Z�0xm$n��W�\���������G��l	�UVN|l�E(��9`�����Cg�H�d��.'7�<J7R|o����+g�~�*���ׂ�-��e9ЬJH�b��R�!��Ǔ�I2�^�C��RK�o��b�蜚��=��gј~@��y�_qg�
d���|Yl�9����z���n�՝qݧ� ��ӷ�1̜�v滝А�YJ�P_�	'ip��G�o�qo�P��蚶:��{#M1Կd/�uG6�}��fQ�����J&�_����rD��%��"d�f�ӣo^,���7�i!}��h���_��F�Rԃ&�V��[�M���nt#���yLfе�d1㖃/�[;�(/0(e
D��|�Fv��V�o�����l���U_൴kq��zF�Z���� ׎C�	ږ����Y��ü�]:�a���[� =��|\���.���'8�mm�h�U���y��`P�Z�{^������6�����;�:H����濪/$J)�+��Hsđ��+��=��3�|^]>:ﵪs�A��7Ϩ~�����N��a�H\U�A;���8�͕��������щ�/X_�j����ٔ:���oNi��A�@��gmt7��"P4���.�jtU�/I��~��+�{_/��K��4]�}e��~��X`���2�o�Q}'$���48��ax��Q8��^ƞt�Vn�50�[@����]U�џz�/���͂{��TB�͹Ǡ��.W�]AZ�8��p�ąLJU���9r�.�r�ii(j��7@'�(��T ��]�2���ǿ'AG�ٺ��Tp�H-Б+̵��呕լ/ͫ9��$��rĆʒjPx��q���Q-���ݹ����]�#�����JK-���x��:���~�OW�e����E�!��NFN��A>�Gm�)I�S����.�zhK}.�ud�j}��گ�����s���1O�1-M�٨#��_f�)c&~���,�ϧ���A�*4b�V�@H�ĩ��@(.katW2q/B��˯�M\�I4z�T�4j6�6.�=��a��!e#X�3����0-�N�~�P�_�D���i��7�^aS���>�R��I��o��JZա��~1K'�o��.}Q���n0W�ee����z�yw��U�<l����SC��#0���j{��ݼ�Z���q�~O��^7����5���t�}5�b��c�@%��uy�4�}�h�o�1���90j��!hc���J8�2���ї��W�Es��G��s�P�xG�[J�U9�Ү�H�'
V^�2�q[�U�l��h4{����$pp2��D;WK�4�J��m>9�~��/�V��XE��7C�hk,S*�M�z�]A%�4�����^�f�1[�}F7���ȇ��}����}�?�}d�s��~���{p�Q�q�-�}�z�AveВ�4�#| ��ӽ�}�o.�ұN�s��Śf�
�O��Vi���Tl�����:q��tS�;�ٔAsa��o�; ;�q�^ �4�h�����9���;5�A�~�$׆���Q@��:bs��Y���ׯW��w�b�-<���������>����<��r���"w�oCx����y���<�2��`�$;	hk���L���:�q���*8��p�LlLo�@�A�8����Ep�Zpl�a����!�A,�]#�Am�ă`C�����='�w��x��8�yZC˜���;L��p��~�1&o����)ov��������0/�<��NB�pQE<V4Ѷj�~m�m�=#�!���h�{��E�2"���A�<n�KW��9�5<��'�ǻQ\M��l���o	��T�ȥ�WiV@��>�?�rT�	�ZP��C2�|�����5�����i�����F)z��V�X��RU�\�tCS��5����\�1&�~e\�d||cF�n�ͻ��)�d�����b8�u�&�n ����5�Ԟ�Q�e�X�!o��$%�ѥ�w�ޑm��Ȍp�����쬓�S�ɸ���||�h�ag���	�v�^N纭�2 ��Q6�令��+l����M��]�v>9�fxz�نChN����\<���?�!0s�z�o��P��L�Ɗ��#���j�9l-���/����)����F_���n߹1���\���i�>s,�ܝ����2̾PFZ��VH�x�8�xT��'2��0�C��Pބ�Y�U���/Or:o�X�����EY����+l��n�~f��I��R�K~yA�Q�(_�֩�h�@���qoCW���i�� kw�K��� 4���O׋Kt���9kO
xo��W(�'2s'q����P��iO<�0R���*E}�WL�e�k;����s�||�uܿ{&A7���.��9O��4��%i<0��
���m������[��a襸j%�K�1��Q�>�PYhcU����ԡ�J!��uW�e7�W�0�;�LՁu��6d�&|i�[�	c�ǌ������x���8>[��]���GkƯw7�c�j+	}f_v6�̯��@�g�_پ�*���V	�� LE��{^�Y�5��Ƴ��mt���^e�Uu�4o����;:�QpÅ������g1�՘4ʢ�ȩ�ҏ�H��m���ҢsT�`ĩ��6�I&�3��+X�l	A�,Hۍ&f���o�Y¯p[�=$E��;����q1��*��Y��3ͻï̝��uF3�'7F+���@O�"�o��;�PsR��ٯ�.�5�:�;`�jq��O�f�\��3A�5R�n���|ś4���g�}`��wZ�.Mɘ�u����*0�pJ�En<����`�o��6��p������SZ8���Zh����8Vo�QXm���:��o)�}�siTB/�K���������Lo�U�\ǎ+�1ѧ��/fM�suo���C�y�Z�)%�}
�fk���WKc���y@�A���m��m���W9[��]}���|R�cuv��ިx5H`��,�|�����h9&\�O4�?��d�/c�,vR�ޫgr��m�����t���a�?{Cꐎw5p�h�+��$Qt�6��1����^PXX�u#=��nx�� �H�)]�O�|�91�J��˗J���U���]�e�?�8X���=��X~��ʮ��F�������������m�XnI�n!,m���Śk8ƺ{��%N�3��7��N�N!��7q�&o�	���6��>%U�����c��gQnh{(�֑�s�aw��q�Xix4��i�{۱����3��_#J.r�N�J��ￒ5wK/^q�ZV<q�A���1��4F��w�xY��I��zy ���n~~�b8�nJl[��k�H�W�[NA��erd+7Q�������4K�n�/=�xV�3mV��Qq�}������
�73��%Ť�ry`J�&������5��S7q���e
��2n�fyN8�4�8x77��ѡ�w�
�6"����|�zR�ⵏ�<�s�+�Q��^�����'|���隵�?X�o&|���YX&��x긃(�<��� ���a���VC}�S{�Ii�yߵ�M�]"J����^�u�v?EA��T��\�$�n����:;���wO���ox\f� p�ڄ��U����e�Ԃx�m���?l����������>���o!�z�R�q�0�T��aUqT�:+N�uQ�f�t�݁��u�Y>=��A�`�]�պ�:#��Ǻw��&�b���RH��0�_�)���q4�1���p ]�}nRޥj>�[��x�K:D�u ��F�H����+\O�!:?�[ȼ�a������J�u�P�Q~�Cc؈�ѱ��gBN���Y)�ڡ.6��QC�UU�V�����i�r�5��{`�!ڌ%����*�������|��v�h��1�͌	�a����`�'٥jF�z�8����g�ui��,���xx��nz/ؠ��Lܰn_�g4��)%X��e�	#��"�Fju#��ŵ���y�]&"������Y��� �r����y��Z�##h�$qss:c�]r�C�f��vMtZj=��Tc4�gxߦO�]9��Yyq�����JI�踡�����&S��mOii	��S[j�Cr��ؠ�Z٦�����b����J��'� �/��>&RD\Fla��R7��O��N�w阰&¦ �3����$�SL1��S��Ix�����q�É|�ˢ��r���n��e��/��XY��/��!�7�jxI[2���a}����)��^{�5�XE�81b��c@y��/�T�s�"[�CI��_�<+
��0�O��&�t��615�d<QF:��md�������p��c�~�3�~u�{yp�u��7��B����]N����H\�n��_���P�}�piBx�8f1�BT'^ac��^Y��i��/(�N��1�1S8�f��vq2�t�S0��2Tx�p�x��R|f9T� {O]Ҭ�m7X���G��;7����v��KJ��
h��\\_!>�b1Oҽ���ZX��6F#�GT�wc�u�ܸ������f�)2|�[�PȞ���_��6����}����c�Io��_ �AI���i�]��&��U��jB�%^�z9��{���m[	Q���h�j/E�2maS��h��F#F�)�.[�qjrg��嶐ܷ,.�K�J�h�8j@�OMz�S�������GC�����.��كc� nP�Fĕ� ��p��'��1M���w��U2�wMK�:g�I��8݇���ǣ�{��}�����*�kX� �s�;=.���|w󣫱ǚ9���R2����!�*�&r�y2���i��
�M.=�D�-+�%u�M�M����k D�O�-��k��"Uʫ��Xp�`�u���ʸ =�q��U-����B�� �Q��\����^������lE|�
b�n ��Ӱ�Jڛ��9�h�Ӑ<�l[��b��k35+6��i�I
����X����G3o��(½q�=��}��s)N9����ު���:}�=��2g���ׯs���ְ��rVoXXح"���垟G�4� ��F��Ep(T�~Q{<�,{@wR��%UA���2n6� ��2FD�n9nw�)��7�,uJb�U�b����ä��"�j�0ʉ��l��v]n�������dgz{i��\�ç�T6�3�v��ґ6�;vT�U�o��_ hD/;m��j��?��^JyV��Wi���*q���Q���j`�g����c�
�Vk9�kv�������Jd����P7l�3���x�놐;�մ�x9B3�"�U���j��ˈ�-&� KOlrҰ���A��T�s��y�<PuϱT��"�櫾;z$ʁ�'�;(��h�Lo��b��#��S��t�U��%a[Y�\�2�A�j�����6-t �vr	9��D�#έJ78��R���܎9���0�K�����f�s�C�J�ѵ�CR-���:�iG�mmn��v*#�7�9��FB95�ћ��př��뵙�K˚8��2�0��չ.*��]elɏ��\x��b��#�%�B�fr+Zg�q�����o���iY�	�!4��z![��§�xL̸ωn��2�%1��2'9�t�,��!�&�I4��7��\������k���EC��qP�]�M\	xǆ"�ګhs_c�1:��X���L�.˗�T����W�ȝt6q�R�So��#�8;m���汑D��g�����Eok�l�m~KS�N�q[xr�f�k�".�cm�;ó5.$������������m��3��d�Dh�TL�?���|�W�d��%���5���8}Fs�mL��@k����O�ҾoW���(�ʵWa`m�;��e
�ћ�{����i�6�p�P�����q{?�/�y�U��f�xgў��O�LD��A�j�M���:U���+�PUIc��8������#�!R΂��cN$S%����M��Did�V��8:����ns�R�xĳ�AT1m?�)x�+�^�C�z��ǡPwh��ǅ���F�9��{?��~�!�d�U�����)��6��p��A�@w�k��u�z�T'J.����k��W;�<�y�]�6�+���~M*/O��|��m��π�����\�2Co�h���:9k!��;�I�V���ou�Q{Sq��|���۰�4pȀ Ug����y)bR�j�:הQ<E�|f2���d7À�z5��Z�a�k��| 7���!���&yN���^��?�t�5}@�ԋ�X�~��"K%���eܧ����2K�Ճ����-�4��0iRxru5��dS^��y����2mG��]���	T<A�������A�3$�����*�]Q����~hcWx-e*aJ�cB.|�.X�F$I�4��]wÊ�xT>5��Y�gMBI~�)����� ��~{	��@�ywz�c�h���:�<a Va�x���������h�M�����+���z]J��O0{��h	�����M>��S� �0���M���X�X�X�u~�C���7^�v�D�-J8������@���)'l��é�w�It1��BmM�8	� ��Q������ZNL|U�U0IEih�Kv6�v��dR��o�{N����ƃk���^��6Sݙd5yD ��v£6O\
�k�M�b�E���.��=�T�R���γ�vD�X ���ɻ��U:T9�ft���h����X��*)�ν��߈�7���}�W�1�>~]{
B�^!,.B��_�*��j�#Ⱥ��ft�2*�����98�M��+�n���uM1J���5�����h��B}�ԍ%5���E�����m-����d/��&�4���*|!�����}�xv���d�R䅮|d��=�
wj�:Č�uQ/�V��1�L�p�� b0o�����G�ݝ������S�q�����YOj����Z��O~�f��|�s����&���;R�^�\*���q.5sZ�~՞''�B���j�6 �quvV�?(0P�s�3�^����]������+>[�j}BZ�3aT���u4-�޷���}�=�X��@>�y�+b_�W�=�[W��L�l����� �r���t=nW�ǐ��_
���͋�F\�aS��u�����̹-���;�G�8K�5e]�N'��
�[��fe�ZJ�6�{ � ���HW���~�}S�G�a��]�v��@͑�����}5�d���,\�/`��A��g��Zn�4yz2�q���Z���T��_�s�ш� ��8���Vb���䕡t��p�̹0�T��f��XU��O羘����<>�:{j"=7��r��ۢU����&A�N��_�Ľ�m����#ǃSlO��=��6�-�/��������g<hl/����ݱ��4���YVh�b)g)�������6�����20qd:�.��Z�J�*qU��o�,Zw�Se;�&�Xn�d*�zL5Uֽ8%+-�q����}��I�κ£4
q�J�8��6��3���f�5-}�{�}ݜ�f_��� :�ϜÐ��"M̍� �<����4�(��?�7��<�o���N�O�(Ȥ^��;2�	+:��c��i�[�=g���*$4g� Rq�M��n;���gu���u�1tK���1H��,+��#�b������nzp�n��Wi��q@	�g����V�������.��/�Xh����[{�H��g����r̭����$0�_���������ub�C)�G�ݟ�^�I���y�\�Ǝ�Pc(<N�Τ�����=Q��`�(���@9�^���}>�K!_�^�PQ��m���k"����ꯃ�*��D��c���\��}�zQ���Sc+�@ �X
�_�1��qk��6���u�oyU��k�tN���~�)��Ѵ��/l��Jʛ�L�D38�,��Zq�r�lE�i���ʱ���\����v�S �,ED����>��sz��°���������>�@�� @��k6�}��2��o!�\�yO��3�Fr6��݇��~ͧi9����_�5�Ɠk=���}���L$��i�Xa�|ݟ:�:��Y�����wֈS��K�1�KBᘓ��.��,��D�D�J��}l�g��'q:�B�Q�	[��� �����y��x:�o��K�5^ۭ�N�h�}1��΍���TQ�歙W\?��s�H���Կ��_p�q[�r#Q܍F���$�u�a�������;�N�f3r�"Ԣ�3����dn��aY�d�3�df��¾�s���Q�e�$��	<��x\�������P�n�N;v6Rfsn<�׾w$/�/]~ xb?	����������8�m�$��������b�N��"uY�vy�3;���� ��Z���G��$�OԦ�AM���(��8�y��e0��槷[dp��w������t������F= ���K�׿��H�o�)k�#o��I��z�}���������O���ei���!���*���ǁ�
� 	�"+�S�)[�Du�=��g6֨U�w[ �S BկR��i�
�����gC4�d���O�p��4�����H�x@�u�o�Q�����p��!��R�t]�L�c�dňG�QP �hL�� �فj��K�z�X�/��|m��3&қ ��qs]櫷o�#<���l����辢{�j18F���	����u��R��M�6Л� ��)K5���˽�q�U<'�ug�;�@K"�\��Q"D�8�~o�kzHH����7S�r���^ �&"�#�c'�H�Ks`�
g��ч�.7ن�.��c����4fP�c�"��GY���b�gU�����ݶ�aI��Ĩ�~ˠp���G�g�1�(�²<Phf�ǹ:>�X�u����H�^�t&���(Y5o� �����}�Sޛ+���7����`iZ�4r�*��}���Ɩ���@!���٧RdhB�BU|��i�#4�m?�ιѤ�4�5fue9��fnK��
�!1������܊��K�>6����X:�ހ�є��vF��q���N��;���(�3r�f>�e��#Efݣ�t
1G�8�6c�%{T(��Jv`i��7�,��39{<흯#}�(��Am�1@�Mz�%]��G3]\*3~����./!��B�>z�֐�% Wg���h����1)�w0N
�Q���n�>����~cE��@�K�|����S ��/�R5�A'T���J.̤������Y'f@��f2eBUy]ӤL��nE�b,�ދR�A<kt�:�WǨ���9���� lU9~���.�Lu�S����	j|G����}��[`죌ټ�QJ�߶N������OZ�1�r��i� ��4�Lplc��Ԍ���6q�'J�ò�	Ks�پj�+˪���=9~k�?�l���J\Oݧ�-���r��f�,�HW8hV�:�R?�����@�� �	�
��T��Q���ؙ0ft�]�~P�F�:Έ�l����  j�B&Ƭn��r��۵|��D���<�6e�4�H�k~�F������H���A��Cv�bx��k=��12���������;�7�p��<�*�Rr�\��ΩNX,�E"A�]�Ӊm�C�Ŵ\�x}ʭ�x�Ֆ/	}-{�noYY�5�����*�l�<c�6gQE�Иy���jTt:g�8~�6^����4���Q:=2\FX���S���$=���]��d��'J�= �,
Fc�}2v_t	쵩�U�Ll��v:H����_pK.([�r�#�0꼔}��Q=�n�=߾u��4T��s5��U~v����dR����/Y�Q��#�ֲ��o;���+��*�>y����	=~��eB^�&��B+��	d��C�W��ǝ��ϒ��!�탼.�����d���S0����w̨[��� �v������ܒ�Q�B�cwȫ���ޤ�֊�#4c��(�FH���el���uG��5[���I��֒D���q�T����Y��z���@�[�G��-�ט��_������=zD �5��*�u�=��8Eǉ��p���M��Db�ۉ������I�)�Le����y�E�64�=8�yJ(��[���۷��IIɤ��C���MV-���������HU�.-�ح&�?�9'8���!�aƎ��eң�yY%��E^��ު.鱾�;;Y���+��q���ٛ0��".�x<a�,�C >��%{�M�?|e��Gɂ�aSܺ���k��<���n��� 7ng跄�G��2������>88oQ�cr�Ҡ&U�p����T�
�.��W�v\�E�T��=wR���ڴ��Zg�)���Wnc��/��<
X��Sc�g���p�[��0�y����T����ը$�K�ߖ�,��?��^ܿ,J߫*�w\6g+�}I
(��@+E�覍��Sd?����r�K
>s�6QN?���q7��Y�5��k)K����T�9?_��>Aq*���^R��˵�CL}�Rm4���@o"y�7� #.K��P��+|~1hŹc�+���&w%���u/�&�� U��8>G)W�����Y�1��_�s%P��˂*q;_{Y�f2E�K�Π��Rw�7+���~Tz����� 嘝����h%S�3s��\�����oS��ũ3h C�;}�a>�_���a,P���íBi���������+�m&B��K�o��.��[�k�8�����4C����ɚ�kL��O4n0�Isݜ0�8nƓ�C[A���A����Ez�g��~|�Z�����}�.@��������G��ƫ(��ᶖ�$x��a���L*��ӿ)(z}d��Pf�����[�y���X{��0� ���:8Q�	��Ѝ��Qc�oY����g�t�r����1U�ַ���f��<8p����� ��8�}v2�|�����]jj�Ǒ���~�O)��<��N�L@��ͮ��מ���`и�����X]��\T���;�?�b���l9� �XB\n�}	�ʇ_����ms���9���J�w�s�7�sss�UTF��U�6�w���Wmw%�ɮ�5��h�I?�c�]в��ge�N�s{��+���{�S��2למSQq,�f��¢�]kkv	#���'}:+�^5��ng}B�Z���cn�8������Y�f�]=�HJ3�Si�	}&��U�&����|�;�܏�n$R������Q���u�������j��	4!���ZKbJ,h�3�6dh��ԯ#�Q�Jk�Tws��S��
�hc�Zq�x�m���=��~���G>�n�L��G�z�y����6Ǿ�s��):���:�����7%E��p���ߙ�ߊ�¥��B	�G���9d��c��Db����;9UJ�7�����3M�y�Jr�N���h�\����-ދˣ��*3����ѝr3����{��C%`�upS���1��)J7��~xe7�X���Gu�����9�D
�ۻdڞ9$������T�H��`b���$����o��������`����>7�15�P�{y@��W�Oxt���� �S��g�����_�)7�����I�{�8��(��";;a��Y�A��ߗ{��q<eJ�/o8=iu7��T���������v������c�7�οMe�qsu[R9MG2d�yB! ��M5�#������v_ �- ����1'��=L��y���[@2���ꍪ��OW(��n�X�8�F��?Jc�of�/2F*cʜ#�+�T���K��M�\��>�|��;����CFK�s�����r��2Պ���~�>'p�E����!Y���ڑJ�W�a��ap*uI��?GС���0��:�8ݲ����љ�c]�8�s@�?��b����P?b rz+���x���B��T�i�~
V�+��m`�x��~�KX�|��DY)�^K�'�tQ�/Ũ��h�����;���T�t(n�A�����c��|��ԫ�x��'���n��+�b�8nM��)����G�<�ỵN������td|9�ΝQ�Lх�29zC���궎�Og��>�>���q<�7���g8��O5	�qY���}������{�)�k<����"s� ������{#�Y�-�`\6���u1=���J����9 E�F�&�d2�_����k�ky	�����b���pt�8��pc�����У��A4�����1U��O�"a��l�����"��Ν��Q ��U{�	q�9�b)�;�����O@��=�.$I�c��,�	�!���0�~%2�J�j�>%��GL�_.֋��G�)�+�hia���s��+$5�ɵ;Z��(���񪮮��ꞈ팃�M�mN��*q��a�K[����8���&B���m�G<l]�33y���z�)ᘚ�$@
���[�ǟ>}z�
#�jp��B�eX���9k�Df��;����"��z��Z1�Y�gf� ���	R����*?�����+����]��P|8� �0)�`[��/vz$�jK�띍�S��궷�$��T�A���J�w2R*�ܭ�-�8�T&P"�
��v:3�4v���契k�w%���*Rv$���b>����U;e|�6������MDmѺf��S痼]W���?����|���;��Q��F����&���b.�}Hr��e+���(+���H-6�y�������jt)�a�1�I�x��Nr����y��r�2�
�l�혉B4j	ӧ�A_9�%}M�8"����b��S�#T���� ,���0B7S��R�K�x���ԥS�m8���/�2�E~���������B5h��oa����\a����`'������:�^{x���@�����f�����L���$�*-�V��'��q^:�y��ϵȠ�E�Κ�!�����6bQ�-%�Z15��aY�ʝ�E�������G��H^�ɫu���u�x����K77 ��U����'�%ee�D�H��ӌc�i��X(e�?$m:z��~�6�g���]�cH"�W"kM6;:N<m�<1�	9�\E!˲���w攵�l��>��|L�&����������sǯqc�3�U���@yU�M���R��t 7�Sn�+Ԥ�J�A_�� �v���`�p��G�	�潽��)��w��IdGk ޿�tgBo��B�$�I}Rl�
��K��$=4�2h���)�u�����][ ���w�\?%eK^#�=�f����댔*�}���\(�v�w��Zdl����O���U�/8�խ6����=�2�&�l]X�����W)%����4K� �Hw*Kw�
+]���*,��tJ���H7�,^���}����3'���߈�zxn	������RC��%c��c��p1�å�Pfط�2�Z��nlB���kT7M&�XY�GFN�J��_a�����k����Ԟ^�r�R6U�{<�&lL6Q����$EqI�#G�Fjv&4�5" �R�ֺ� ��!.���J�\X�������fN\���:R�(��C��L2��r#�tc���,466��~�}o�4޸�ox��sXo���P�3`$� O��<���]y���&�A�!H����[_A������8���x�Z�� #K]',���e'����o�kZC��ZJ�٘�w8����f��®��f�fYM�S���K���7����yծvF�C2J3����E%>��Wc+Y��h��>�Va��耡&���7�����b�R�1ӱ+ �R�>s�pP&���Pr�DX�h�<q�y0x��LNrW��v_CV	�_M�^*)(��bk{&����V|$����:�{K����:��屄��7�uҔ8^Cϭ碓�	�b��[)`|!A���g}�����^�F�����^��w�v�H�sK�+��z��ǭ��@;�D��|YWW���Ij���T�����	�[���sc����V�����;�׾ڵ����=��Έ�x.=��3P��O���WG<����?ZY��E�S�!��؏�O�!]O^nQ�:��D��^Y]]=L��T���_�܆���L�0���F��٢���(�L
m���K��>5�j�b�i��(UV�$m�k�����Z8Ԕ5�#+��l�.Nqv���DU�bSn���a�%�����`:v�����5;	�����(�6����'�}�nY��;��컩N����~I�~�T��4i-������ȉ
��W������	�S������>�4~>��:�g��:��˵i�29�"έ�R\4�#��dش�D����)��S��V��fO9�L����}�3r7�2w��Ja����yY�`z�\l�����m��4	AS���Ttj:+=|�M�R̡2���k���ķ׶�X���LoG�Ȉ^`��T	���Z�o������]�ñ���ӞG]����W  ����_Ѥ��W��^�J?����*���7NS�[%�]�\��D��;5;V#
bꪜ�~�(�S���R��~%�(�t��V��[�L����co@[k�J[��Qcf��3�s��R���=^��ՐW/^��/ԇ�įL�:���9[��X��-z�T`��Q��4�F�B��/
u�
�D̳@?C˜� �ٻ�D�$�E�r��(��R'�r^����sE ڪ��G*Q��۷�#
a�2�)��Z�����(^`��鿴�
���Tttt�s	e��å��W��i�IFbA��m��������N��獆�=�fg�:y��T�����hh����s�]翥���=ޮ����7���.����}d����y����r���z˗���K>	�~ީN{ppP`�:g�z�@�oB_9[j5x%U��	��J'˟�X?_���e�:2VN�}����ff����^��W������#�W �1G�����r�:a��b��#p˽Mlp��o�;�}�r=�#(H	B$i������
�ߺ�;�������e`
�?��L2Ͼ�!�/�:t������V�4NNN��&���R�A��\��$�PL�x��Tc�����`�>O��7_N�GU�*(�323�����\����_����_��5�oJ]CCԹ��]##�`�����W���S�f�o���)o�h��-��H]"�+��KH�?�u޵�������O�����]cc����]==��^����NLL�/�W��X��t��EhtDDD���u[�薌����2����+qqq�[[Ҁ�⿅0Qd*{l.����GI����}�
hxf5Rnׂ��u���f�ꎾ���֦��`]}}��/�r	(IeeB�Ô�l����􎯒����ߔ�x +ۚR����{���߂
o�����7˱B6A}}}fffQ!{�Ći�X��Z�چ?&�
$�q��&;��Y�ntt���b�W�`2�6775*������%����gZ4���F+vww�ݑo�� �vS�xp���qR�S�����-3��3������&��g�A �B����M��/t���|]�i5�qN�}8������H�� lH�Gh�ߛ7�������#X�9:�oni����(�Q8�6�=�㷌�o �P�o��Fi~�h��_�ffi�.9bт�z���m�V���Xn��� 8oB_�Gh����Է�����jr�r/��74J����-����cNɩE�G�n��ۛ��$\^�[C�O�Tݗ ���p�wy�4L�1��S�t���IX�^���.����{�/[�6ek$������rh��$m��?.��Hȸ�fB<c�"j=: )��AIii�S?:J��կcZ�x�	e&#���áW-�C�����〹�ir5�<�$$�ہ������
3��k�!�o�8�̓BϝU���C��-��<k � Ov��vyɃ��X��H�4P,�}�?�����7xs���������ۧc�������������i���x���%bb�u��%E�H��J'E�[��h^룗�:chsʯ�T*Ǌ̗���b��D�z��R�XT&D��@8`�L����-###��Q� �%z����}�����	��;uA �Kz��g%�*Qdgw&����!@��1����OEE|@a���9�؞O�q �,�۔z(�\�/�*��l.�I�U�m�ID/yt;�*��}٘*���ݧ��D7��od��y���N��G���������ʆ����o�F��w�H�j8dbBmLf7<�v�8��j�t�[B�5ZZu�H˽9������P�I�?�.�y� ��0*̀'chH};��p�HrW�f��`����v��V&��az�w[_u���<l�������ͧ6����\\�J%}�C1�����?��l��*�un-:���1
?�x���

�4C�hK��x�.��<,�uI#�k��b�A������.=�zooo������GW� ���l����U:e?+���;�+�Y������ �L�%��n}'1�����oݒ���ѿ�h��S�$�PE�R�֎E�Π�x+6dzkOUI���C*}���㑮�UXXXn+6h"�RaZ�	)W��9���4=ʮظ�2����B��CqBO�(���x��{���->����"���%%��F������ �+
]�	��Y\��x��h�_���n�=�� ��d��*-��o��H@�W�$��͸�쌌&����z������]r?9T���{�T%L�l�CP�0��\��kk9;�g�?�)��}�S�Y�!ƚi�W'f���x3N��6�J�ffgˊ���-�6�8˰�'�x��4��x�}LM�.�~^��CD�TVV�H�7���^߻{���K7~��L��xv���R�Vjʮ���5�I~ܧ@��a]ʿN<�ƞ���N�M6�U^��j�E��z����x1-�mKK*���[��G��	�'5�G_[JW=co�g�קv���6<k�m<<��=<t��$�\�ӹ~7���CU�x���D�8���1P�D����͇���><s�Lޒ|Ł�&}��#���n�e�S���@���R�VS�Q�L9l�P���b����~�k������F�C�v�I]���������z�[�Te��˩����� �9ؠ���z���d��0X.SfQ��Ж3�4@��LW�(0��p�4@�n�Ȍ�	���w�g�d�Cz���!��.R6MM<թ����OQ1X�m9�K�D?�Gn�����dQ�搛�;ۋ�<�뛛�����e�X���� ������vv��\e���@TLll�#&�3u_����H-�?����~���x(s��H�u�J_�OC��|��������d�*h\,lJ8/��w��g�a�w���V��nu'q5�g��d�����b����� 7������֞�(a]6���]]�7�3&/󱜾�F⧹d���-����b�歆� ��Z�>>1���0&�$���
|zck�ʝD���W�V��.ՙ��3AH��OE�-))	I��x�ߑ��.�V����Yck>�600��^�u8����5y)�?��	�����"���]A�������������𤨇��z�]>�c�27WNc��=wj���Q��>NU�ߖ��m���L�C�����8w��͎���lK��䓳<j1�Y�㣦�r�AMC���X���amY�eTTD� ���g���1bf�.���8	�������y	�O��z��d:Q�R�5�Г��E~z��7h��M6�@@� �V ����|��n�ؗ���sf>=���Y�^C&�C�%��W��*7d؉��K�ى^������S�[R�XpD+��?�K����<M��9����@�Y�)�L����������Mv��F�G`�c���:�z'c�s�tR�i��ữc���w�"T�Y��Y+5�vq|$�uư��}䜋�@W����{�������:��#����BBB�yyO�g����9���g ��2�I�S:�P��ǹ�睊�c���Ǟ�ǯ!^��_���V�Xՠ�Tˬ-~�!�yyT�U.��¿X1��H]S�j�r�y�W=��B4(yyٚ���r�ڍ��-���ytؓ�P� vl��4��c?�
|�D+?����(�d�LI�Ǜ�E�/V?�R��!��=�����}��h�8>��tP%|�x;��7�"��7AЅ���/�T���.�8I: ��E��$OB,��ؙ�lZi���1��k����F��Wx5,HHcz����jd���f	�����Up�0�w�n� 8���dE��2

���쇚��BDEá́�O3�u�.��ﮜ������F��tp�p�X����f&��|4�%�ij
��0fw�x4�]h��8���/A!d���~� �DMQ�r�Y����`����i+%v����u��d�q	љ���s�f��-:���:�[�?̥�@jME����"�b�е���w�#.{r����?��J>>�.I���P�q~��������yw�?����5!&;���^5\z��X
t��G�J �?\u899�99U�o���߷taqQ�����.���I�1�����;�p+�T�M��օkྼ׌�������d__�5:��� ����@)�@)U-�,��@����Ja��YUUî�I'q
���F�Y��߸;+uP�G�)����M1��/N��˷�.4��Ns�w���@�'�=e���=��٣�{��V�<C�k�c;��؎j(K�04a7![@�R ��Y�	�J-�'��S���A��_����ZX^Vc�Mg��c{���*9��aq��j�@,m�M+�����1q����hp��n�^�� Hmm����rsU��31���0�ZXl�j���E����ϯ-���d�b��ъ���[�ŝ�,N!������R��C6�.  O
ZZkFC(�5x�Ull ��b��^�g I���C�b<�v��ٔ!�2ꦎ��"i !���I�� �4 �Aa�?Tb�;:�k%h	�b��Jl�3V�?�v�3>���e�q����.شւ$�m����D����!# ���1g+��7Sɢ� �d>��Θ��ɫ�3I$��c�T5�RE�u���	5���x ��[M��uT�m2�� ���R�x��V�(e��ڌ�<TUWϮ��JThr�hS4����xg����|���I�~�r��P�MB�����Z���+�v�R���� ʚo�Y�^qԲAU�iƚ�}���q#�C6c�XQ�舾'l5����� ���t��̥O���n��@t:�	����OJ�̴4)�����W���j���k�dl�����-��s�v��EH#%��
��Е�)a-�`���X6�i�-�u��z���kHb$�PH�hm��5kcl�����Z7zp��<R~8:�����H���)�^$��`����:����*qZT���q�23�1QO+�s���9��I0}<�X�[�x5��*swn��mw��j�W藉9 7`��^������%�^�n��G�~�9/�h��|"��<�*���N�%Tf�A��.�ӷ�N���G�EC?^h6)Z���B�~������x�N.��եH|钙��0KZ	�ĵ�N\��#倇�O4�jw���z�0wuIۢ��m������	wK3��d��� ��r�s��j�U�&'i��VB��=}����y����q��=������a�v��ʘ�(>|���lUs��| �����ѭ��B^UUՓ�n�R<ğŧ�)���a�f@�ݜϢ 7�>{�yT��f�w"��}6�g?�r��A��+~��C���L���~�:�
+���;7w��J>�UyR8�YA� ��Ԡ�ߌl� =\zm�S��r�N������~Ȥ��6}I^z4�֡���U�*��h�!d�r3q|>�t�K~/�Cl���1c(�塿������@�[~^�ey?WFwUdDD@n ��N�MM8V�O���++�zaCG�^^5��H��?�(�}�Ձd�v��+l�Gf���:���u�i1^��g ��6�Nɤ��Z��B�D�خ��5Ͻ��ƫٴ���FYY�B��Ѣ� q���b�ٽ�Q]�s��M��ސQ���B����g��(l��2��:N.C�^=N�c/P��Y��Q�BN�{U�q�PìA,���q�2}�@��HT
B_KT=�D~��?�����;p�i؄p4�=��D�� A�Id�{�����z����A��J�J�c�5Em�V��H����פ���Y�B���Th!=w���ڽ��CV��,zw�_Q�����J��ڠ|������KY�Ŏs_�<M�7%�\��k�`�����Δahxr�(��?�8��r�?�`���W�S]H:����t��()Q��a�G��Q[����U�\Ba��ҹ=[����w��a޾�[4.��|� (���:
= �~�;V$/ۻ�]���Jw��Lށ��jjF���(�ԅ?�vE�� �Y��G�`vYp��(.�wk�M	��;����P����mL��o7�E%���6X
�(M-qXm��?rwj�๪"L��F	�^�9��C)��+�V��ҁ������ggg�J����E�~!~c���.QkO�\���}ZՈ��Z��\hh�V�2�}��~�P��M�W]�pK@�ٚؖmXb����@)�ԹN�ӧ@;�����}v�7��b"�����iI�#��Q;Z�e)<�8�Q۟zn\��/:���gk���6y�l�֋�$9��TB�-�U���.cOY�m	�O��j�IUE����^�.�_g��:;��3�k��7�j�Xk�I����P�#����Є�3-	�W�?�G��s����e�U�_�!z�\�RT��;��GS/	;}p���4�N��q1�YUg�r�����������wc;�fz��\��*������m5��q�l��������	���9� �K/�	=[-�m�RҾ�Ψ��B��U��W}��E$zGΝ�\,gV�Y�y����&��t��&����� �V'�	ș����v=����b�ϋ0T���Q�;�Ui}+��YݵCqRg�K
��&	�Y�^�9�]�s�Ǆv����H&��`�"w�kV)f�� ԅ5�j����,W��WP��Wt	���N=����˷�m���b�g�+��f�|�t���r��(��aƸ�O��v��ѝj�;81|�
gB}������ùSV#�-vL�AW�ծ���f�,Uj��`�%����7�A�r��JE6�N�P�LEk�𪟡f�T��L��,A�d��5¥p���z��^�2DnիM!�2O�%J�=8˙͛��H+㎗����[�1
���;��5����R><1��}G0����(�/	�+AT���>=�����s�B�����lf���fw/n:�\#9���-m���PZ�9���¹��%e�qf=�J w����C_v�S�;��k��
�i2�Y&K9wfګ��o�Չ?��E8�n��?θ����ֿ<�M�ƙ'��A
s�Ke����9�գ�ͰF>�<W0a���n�����5ˍD����!�=�7��}4x��Â�]77^�.��ݚ,5-��z�Ie��}:"���)�,S�A��biQ�T���oD��˹�b܋gp\i�6��}���&�U���X%�٫����L���B|]��fK��R���Ɖo)�1jѲw��<��\�s��w����o���v+f�1J�e��!3���[���b�A#gv��D	��(�� g�2�$/~�r,��U����e�sAS���QA��STXԧ�\_���I�^�bկD��K�F���K�W�?�
b����k�y3���j�z�~\�A���>1��ה���vl��ӭP�U`�B�2s�8��GLӶd�<7���S������L<�.�P�9`4��P��wd"(" ���!��2�Bh��~�����i�ͩ��Su�Aa�2�7FB:�| I���̰������"�l"Wl����]��9�:���rڄ�r�Y��J�ƙ!!��g��z~/D}}'70oC�)*e�;*eK���|x����O`���w����s:.f�K��+�ul�p�i�c��zu�6�}��O�td#h����+|ٗ~X%��d+9��mG�����T��B�J�� H��]��/�b�X�]���`�v�=�,���t	ۈ�LM��rC�i�}oʟU��d+�hs<{�Ԙ���R�mP��aZ�v�\�����j�z�Lq�!�	@���T£�fn!۸1��G���zr� }��_���s�rV�>5%!��ک����w�{{f��W��H(s�w��$����E��p��'��d"8rY��S{�����\G)��{�PKE;%�1���.*�<��!�����/)<�A>��!�ckd-�+�슱������m���*--?�N7P`ZXY�ӝ!+.5L~C&V�;%��:*�Uqf�a� W	V�fiQ�@��jB��U���H:2�����Γ5��1�V;W��*����	�;��p+��/_�����;G�#&�·���#z2�o�{���&��ϡ9T��¢ڣdE��*�v���KUّa�#Di�KRj7h),�5b���N��j�o��e3Rj�<ZM�\��勫��#��Yw9麳�.]��0��~��:�����!b�z�"l��"0g��Kɔ5�9̻��,w0dw�c���3V��߿�L�^�b�0Z8�	=�yJWW7�������N�Q���så�s=�gL~g�Ɍξ��t�����D}����kS�w76@�*en�%`�	x�3��GX�:i�AӾw��Ҝ��4��f����ہAA1 o�Qv=��0���{����l�=�F��55�����!q�g_10��-MwS����"?*��B(�i_�g��?�RS���yS�u��Nh+�۵��S}cX]ɠ6�i�#�(sr�P��tHt�/o�3Vā�4i��U�Wk��r�W`����T����g��z\�&��� C��UQLG�Uo
8�TK4�I��aٸ��b�����C�|�2ā�C�{s�@N�=��P�;�k5z/Nu4�-�?Si���W�C�f�r�"ʝH�z%�?[F��;ܖ9�d�U����  �}�|U�ec4�;}s��NҜRj3n9����x�A�I^�v�kI߫gyb|�BG�yI��if�ߍ�)ֿ
�E��teRl�����s���f��
�ْJ�S1*]:��{.Tk�O��E�ͱ�]��Ra��M�X��v0����zd#�-�������R����밴�_6�P�^�����InN���6�����k_��N%~�d�2�HN�MʦH��MW��M��.c�\�(	�2�;��9�-?�4��7?��a=�(*R�#����\��aܓ� �o��9����m�[☠_��=<���D��)��z8��p��~���Cyi]Na��$��MLM��⭤W���}C�mq�����MrC߆�\Ŭ!O��k���	��#�Сr;Fy(�W;ڒ�Ld�(�PP��{�e�	)��Iȉ�~ۏ���@E���[��TfH�������2:NOXƄs�}�8s�w���l�H�C}��9,u�����yi�)伂-�(�	��z|� ���*���e�t0����d�����5���4p>_;����c�U~�P�)N�떋[��q��*�m�v0������ϋ	���p/���2kk5~j�t���ͬ�"��O �JJT�+Ia/>����MI�WN����˵@Ft~i��q�Q'o�OM����8�u���p�SւA���ͱ���?.(��;�3���l�����U��Q��t.������<�+�ic�ذ��VVPNNN����n"����7��|mn�����[��Ťʝ �ாL SM.�oƩi"�����P�)��x�8����gપ)m��;�H�*9���ҍ�v��3�����0�%Ҩ�<=��W��Н�;z�t��c�r�D ���v����+��-���[}�
�P��Pf_4����|	���ܷ"]!�ޕ��@��\����%��<s�,�܎�fFb�J��2�cu|�� u�\�vY��9~� ��򟾜�Q�[U
��V��Y���c�,�q[��ݜ�vl��I�1�:��y�Ң�U՗S��z�b��W�|K��v �>!�)h9�l:Bb����Z�U���|,�p?�'�_��Mp`#)d̸��Gz�4XUR +�wC]`2%�������"A��+�eJ�x�;9:��?��Va�r���,��B^*�����"�;?*,ꉱ�v$�ѭ�7�M�h�D��bh��L�޵s�zSh�2y�~�ah�CK:K�n#)�~3nͭxǋ��>?o�;��(g��u9gx���-���	y��j��$�iiR�{i��FJgΜ���B����Უ��ot��>|������Y�I��#��GLL<�1`���dIKro������Zsq�����1&��͟���IM�AV�ep9���oN=�F&8�V��K�̖��v5�v��yl�Q���%xOgk)��3-��,�Xٱ]6�gZ,���Ιm�]�W+���.�)���?��UURJJJ���b釫Nrr25H$Q�G��S�Դ�=߿:�ܷ��EEK+��g9��nL���� ���b	1�[;�D���aUar�7�����-ReIW��-I����Y[�|�p�s�sA�E���R�-�Ĭ�F�8I|�S�G������x�>N�pd=�|�&!�$f��M�]���V9�r��k��!c�[�Nk�l����Wr����S�uvz�}�+�*��w�Pl{�-6U��f���+�	�T�Skk%666dB����'��W0]1�����RH6V��P�5q\I��z���|�F�\�����_��I��>R�X�"��Dr,�`�/B�����Zq&���F��`�˵+��i���ؐ���I���/���NS��-?�GgCϣ�7�K�e�������8�z%�9O.�,�а��C��@��4W��5Q}�7�rk� #�@;�y��_�A��+!oYx�j������gg/�7�s��ue�	LF?���vL�誫ke�!W���F�K*l�d1�_<\|ҭE���y����A�{�����H^��@��'li�S�{�t� M�F�{���+�/T&6 ���:V@0�/1���IݬdO��k���� �'�'�/�^-%�q�s?�����J�=�����xWT���g]����YV�������a��6�����A�b������#M�Z_	�c4�!X�.�U�)�M���)�%#=g��y�ˠ?Z8qȪ�o�l���0|즗��.��J=k��{�7����~n�Qr�5)sɹ��g�U~����0�VlN8��m�X�Vb~m1���謸��0���r��~N_��tj��&а5?��{�)���*����%^�&y���	�ڤ�z�WJV��%�s�����o\X�ٻ(�
$:��Nhfrˊ���vB��w��I�VU�zx햍��nH�5��+C�շU��Uc�����Z�]��$��<\&\"Y�h���Q���9�2�󬮎9R�aRI�=x
��c�]�-"_�q1G���ʻԮ�O=��)��#�	R�)�*�-mU�1c����07k�T���⥒$�o�M$��պ�)?3b>�?U�c)���W+{T��L L�?��}�Arşrr����,�����6S�{kHG�u�����<���7QT��	�r��(t�x@c�.��6mQb�������Cc{'[mB�A�pHs�J�G����ZӝpF̹��U"b8��b�I�x��s�T]��0�|u�<n.z~�+ɂ�H�
[��c�����t�
-^ڷ��I=���RW��/	��3��h�n_u}ǁ@}a��a��1_S�{�%V	�>�^KꤿV�x7$�KM��]#���#S˄j�üeHs�s�˪�� �&+�B��N��d�;��)�Ls�Z�ݺ������g}�����&ӻ�ɠ�d[�Ļ8hO^�h�]	Z����!�Q�4�� ,7��s��h��P]kԷ�10����I��y`j#��9�r`�,��t�7��u��Pތ�ҺV�����#�@-b&!~���йoY>���t�U��vp����\��G�jv)�Z[a��z��DI��=����hT٧!V�k5}������o���>�3]�[d�R���qǢ����H��!�c�քKb��t]K�V�:��`������X�U�1���T� ������"�+�=#��ڌl��䳧<a��Y�^����A�-����ړ�E�a�}�Ӛ�����%u����ݚ���Wo�#wEyN�[�a��7��]�l!%�<���b��TZb�#���o�.y�E�+�.~��D�Sd�d��O'vY1W���_mIa���	��T%8�U+#��'.#�F��2D�U_A >�4�9	������rh�\����2vZ{o�4�I�U��G0�p ���RHʄ+4�VFi�A��ha͵�s;idFZ��1��Z�e�v�q���1?}��x+�!����}����~JUo� ;'B��~H�?XH��x��pJ�=D�!䍢�h�h0Ԛ��ƶɹx��!+�ƚ�%wtS%p�u��ϿU+!�J|��튍���������������tMa���KZ���}40�=j�����%9h*�x[:c��A��d/G1=/�RZu��YBݞ�,`P��s����� .���98�^=KP��H7�C�_T�

	����Y9��7��Q��<ߗ>>H�ֻ}�ұ�ʹ����A=���2A���>��e�:�xt��Ѕ�8M���D���b-�����ț#�M�&&ٗw�ᔼ��5��,��H���}�I������s[�f�e��Q�|�*��;�6�;6���	Y�ܒn�D��;�
+�
��х��.V�}v���0w�>�Z���RN����p��2o}��+��ǯ���$Ӓǧ8x�e�-42^�-��N�9�V)�����s>^5ǆvk"�yz�k�]xoq1q�1���O�n�>��g�J������Du���$$WD�E�5&7<��5�����Q�����V�.�s�й��h���h���~�T�흣�j�ru�e��;�������ZD� �a��Gs��NG�鿖?l{;�$Q����#Ӓ:T;덾��Q��-��LQ�����c����	+���LI�a9V؂��+�;���>�C�vc�Z����~4d�8)N������������=��)�d�8���0jC�M�?^��+�ן��f�U���.��"%�I��QoYi���go�
:7H��뾻
I�����Zl�� �oJx׺����K��X��rg�UU_�Ғ�>���@(�?B�2��k:��B$?G�\�6�+���ь�>�N�P�c��ƃ�;Gpޠ#�ʵ��B��T-��>Ii%�����^�"I���=]u\�Ú�ƞK��,^cq������6�v%3H�2�i݇nZ��!��DK���]j���^A��ъ&����(���CV�����e��U���E*˻<V��[��}����]n[:%-����>n��E����$�&!���8�x>>1~���:���ײ�צּ|v�m�;�F�s�G!Y�A��o�m�gnX�h		n~�XJ�@:���n#���,�����~��ò�W��:~ó�ٔ�~'������g���Q��>9�/GӦN���ZWn&|��F�\��|�Ԃ�sT�T�2����KI����������K���B��
K���:�wf������;]�d�8Uai��(ϸ2+�w�nϻ��/�fCM�e���W[f�8w�fZ4�l1K#&t�S�v����2�^�59�
�0����ܱ�Te%1A'�T��e��8�M)���p�f��i訚ʪ��3f��n&��͘oy�!G�����g����T󦝇�myD"���"7��:ڻ��q¸�A[�0��dd��
���P��e;�Z�*��T�pC�f̓y}���A�M,`�D*��s��!=�%�A�<��c�O��1�Ru(�5�����'���*J�й�MB�>��3Δ�B�f�%|,i�PR_Q��9��sY�NǵG鎋�_����he��B���H���>̤zw�����+V��(��i�Ӻ��2�Ў�۽�zp�GV^�T����)��!��іS�,x�1E�j@ߚ�	�I���ß<�.X�����u�RvYx�ɤc<��۸D��QY��N㼆3���ÕlY��
�t�{p\܉���#K0��kL��
�n���17Ar�ҹ�Z.���'/77#M�����aʴ=ެɦ���_p�+���m���k�c��t˭�����=�������F���8� �t@�O1��te�
�#83|B��څJǄu$�����
j�eX��U)�s�1m�4����ؚ]�E��|p����:�U�,��X�氞j�U�K'������+ʎ���?�6�0'���	�=��1��Zm�x����8Q0��,@��AEo�癲u��@>���w�N�������7x��U�1�K�Έ��x�c��w�>g1e���r[���cȎ1�4r�t�u��$P.���Z�%����e�>!�s%������G�-���珛ch�}Q���m�
�i+�b��XX�B���a�i��l�oz;��,�_S��"�9���F�,jk�'�]0��f���n������ۨ'�+_�b6�̚����򼯠cYv�G�޼U��2�x[H�!�Axb�U͈<+�4"ĸc�n��k��0z����+�,��F�r$��	z_R��x�_�v;-a�i�3�I|MN(nn�Ĵ^7D�E��õSU!o��G��&>Ω�MN5�N��jkЛ�B�ý[���ˉ��iEK�Θ��O�r��T���嬅9V����y���HQ�C!D�o��^��W�?d�IM|����
��
�| Ʉ
f�=��$�_xG���Xƿ��$�&V�R�_L�b;�܉	�8�����	F�Ɛpb�B"��!Y�y�X��&O��}� ����8�G��u���Y�sn�Ee���	ۅ���tzmr�Q��(i�%}m�EoV��b ��yE�s ���so�������|��:����!]�4�l��'�KA	�:�n�3޹��R���h"�>��آ���u��k��,�zn�1 Ly�WF=��]#X��!�>Y 5��̓d��ˀƯLI*�T�Y/����T��a�\�q���6��hcI�x���=�X������Ԣ7� ��`���j��Obe�h)C����yQ�����������r�?�!7#*�U��_��v~�GA1�jm:��(�ꐾ�ߋ R[�Rk���pSLQy���Y�����uƋ�ܓѬ�Hp��d�8�bp�r������N��-�c�2H�g��(�]+|���&���d�H'T}T�U�۫w�����;A��_ԡw+�VUʺ�I��_�a��t�,�g�vDӪ��9ͧRF ���([��"�s-�k����;w�P:e�@L�x�B/'����o��3hn�,�IG�Kv;���H]ĶP"��ˬ�	ե�O{S&�	��3��ä]�:��	�����+ɭ������7Nl�����f������.�������2��z�1D�����ѻ��/D8�t��>�~ٞ-ɠY����B8�]�`�LxP9v0�9G�[���:��~JowO��'ٴ]jk7΁,ș��q(�~Ё��z�O��q��%�ڃ=�x�'N҉��%��$y'�k�T!(���_�V��g�)�r�.D@�GMգHk7�Y\�+w�)8��Q�/RUq!�<�i�N��Vu1�BLD�����_-$��F<ΝP�.ྑ�t�ցT}Tqޢ��L]����K�a��7��q�>!�6;*eF���7nF��=h�_z�U%���u�}�d�n``�Ҩ�<5���jB�u�j���|�E����"/MȮ�bd�(�"k�����|l�Rb{Q�����%K��p��[�G�H��n27[�����I!7�Zo��G�L�LI��B\$��l������������T�!�$���E���FXFG�#m�x8T�o[C�I�@c�\x?:y�C��Xf�M2����YN�cO��^N��3.�a=C�C�K������!���Tm��j��ô9���\��ڒi��匔>�s:���ºw��R`d��4//WL�^ʴf�_�Cz��]hD*� ���ԕ��<%��4ܿ	7���W�6���������K��}S�y�^���܋��<=�N����*o�(N��U�Ҍ�K?��x�s�|{l"4K4��u��W�א%j�p����v�`R�J�R�>=@#�j�^0cɡෙ\ωs�ߔ�
��gV&LD��zS�TG�����������t����\�f��N=�����1�$�=_)H=�Wyf&�uS
�l~�hl3s�lh�砾B�iq��H��,� ��q$
Ő���/��*�,��$[���?�Ye��z���Hܜ%z�{�5ө�i"�$ktYV�Fg��O�T��Oz�M�g߹nBF��<4�{v�z�p�"���u��>�5	��8e0��1_��n2gO�AZ,���̽{�<cI9Vi�@�?�B�b�75�ߧ[v������Aqu[ yyn�IB�wx܃;��� �K��A�C#�K�	��xc�6�����n���3?曚�*���k�g/y�>{sJ���u�%+��%��$��_��-薃���e�N[�S�<��
��W�����͓"(�^p�Kʨ�_���+�S#�Dth�'eH��R������c_]7O�-T`�ޓ�|{�ApW=gØx�M�~�ș��ϧ��Qq7�W�����0�>9�8`�П�y��qǴ6�\yG��DA9^��<��.�|�}"*|Y�y:�
���N���G`�k�-ז�:�7�����qk+�*��y����v���ߍ�d���"�{AY������8�j�o��W�i�ى<%����5�хE�À@�o,|ƍZg�ҢQ(FtkU��7�}%0�����aŌ�dwz�!���8��Z
�����q'D��A�:�Ur��IX��J�V���|Ɗ�;6 �I�{r 
V�j�!/��5�n��-�QQ��E�1�J~Qg�D�q�ҏ��ܲ��N��sƃW�� ���ǈb��X�e���r�c��(��C�u�w�O2���R�����L6�O��_yݴh� g$n=v�����U-]�>��M���}����u�- %�)x��ţ�u�� ^�L �zp�]��5ʛի��JH�]�j����@��ӖR��o W$}���>�;^5�A�ԏOa��j`!�-��]7��`4�b�F��B!�NG�{��n���@^�Q��Mf�Y�?w(A�d7s��fFšÅ������G��ͭ�|���~�ޑ}@��J��8��z*�e�R��'w�Z���⋱XJ�	�����-��wG��< )#�zzjmg*�?�{L��r����!��\}-Dj�­�w*�����]>U�0/X�`I��3���&�ua�xIa�C��o�v���<�(S5��9�?�.�t��U,;^$�΁�
�V�N��R��W����F��j�Ϥ*xQ��|)��N��?�#*��[4.2ɏB�m�Zt8�o
�<����W2�q���xIj�/�U��gK�X�,r ��JM����:K��4�F��7�q���}!M� "`SE�֗1PA`pCE���>�+m��s�#*�2~��ݲ	�|���}��3^��
8���`�p�����(|�C j6�O��c�!���Xa�+	���^�mU��q�c��l�6>�������x�Z�+����y�A���'JZ��ҭ{㌇�+��5�,��Y�֥��\��I��m�]_Fr�%��7 �a!<E�x�d>s;!�31��r�<�h�;�=Z柨
~���n�X��ٺ��*���p�;_ngp|_eZ�V���az�6ؠ�)�J����۶��+C{P��o� y0�h�� ����3#�t8�� ���͈ �]BP*Ͽ�s*E��]��xU�L`4�D�r�@�ԏ���A�l����G�K��'q�n>��]o�r�Pۡ��B	7��Wv(�s��;Om�ݏ+�8˫�%�@7p�}p� 4�����m�^�����?4�*�e���ϕ0����yp%����C���g�k�^ފ�8
�WAOĤ��u��QP���� ��  H�dJ�W!�_Bc�����k�'��c���q�+i$2�M黁f'�f����.֢��	��cݼ��qw5!F3jd/�����R�	����^�������E>a`��D���a %ۛ3�ͩ��'{]��~����fSC��Xʴ��%U�;�Z�}tل9n~n{���g�?obz;]-� �I�`�ڸ���<����8s����Ź�g�܄AY��_������!R�@j�b5���gK��
{�	Eof���a!�-�_K�Q.�r���gTUq���Y�lZj��	����UyhxޫwU�T��?�XV�#g�8<�v+��̆_�!�K�W�y'o&8t�T��?��	#�TK��q�Hg	�ɺ'B��)G���?}>42N9� ��� �3��OĀ��b���@���<�9r��t����oIsŞo���11��fW�ޞ:���\��}[�A���˟JR=,Prw���ӯ��}@�0QN����2���Ty��1vO�ط����!���H����<r�:[{�քe���2���z�eʣuS˶*H��/>+'�_bKU����X�?q�M�lH�̍-'�� z<G���Z��c��`�ʳ[�N^����r3	 ���L���Pr��Bd7���|)ױH�O*q�U��z�-?�o�y0���^K&��Mw0�� qe3]�foF�*L�|�*�b�Aըz}��̞� *O����m䝜(O'�iMƩ��Hʛݥ��%���WP2�T��jb��T��`[7�\$�b����Qw��Ѓ���V��%2�f��e��3��]T�}��W�D%���f���S��MH��M�ȆZ�&�����{�s^�cP�\ɖaV�pސ�Xh`gS�����M�]��N�ne "�D��PQ���&�O��-�B���ZN<��MB�ܲ*ß�#�v�X( ��F�e�>�|7�3��0鍽[����0 ��<��S��9P�v��ă0�/��l��w�ܽ�9��+9>��z ]�N6c�L~��W�K�FZ��xZ�|���G���=��������1&{����˔�_�1��<�w5��=�N9:�u�W�r(hc�8�T3��������Im�&�-�U��?�M� �U\A��� �cË�Mgy���8� �t����͟�#����?Ӗf��C��<��`�a��9q��z*���ê�eߏʀ3�q:$*���W`�4�{n��V?��\�e��t�(׎to�����Ɏ�_���ϖ��QEA��� �w���F7ƚA�N����}�Ӌ\���R�����q���Z�>�
���\ȣ��3,m�y��ʁ�U��6�w�����e����/��j�}`�+�q�ȷ�zi�އ@m��w� br���z$������"e���?̻������R;�#��=��ɏ����˫<�u$���AY��U'pa�`��u�}�;rb���N��x(��-��QϠ"s��d�]����Sg�	7�'���q{���	��rT�2�5%սx�Σ�Ev��[29��``PtK������ٞ���b&��*�%��Z��&��!�����`��tQ�� ��l ��m�����9<qD��g�����;�G�ؕ���̻�j�Mj����C~��u �����:����(㓧�b���p�ݬ��R�ͺ�պ:��2K��}@�)����5�&a��b�+�z{��v���	�S.s3���ܜ����}��j����syA@��=��<-�=�@��y95�;�
�ïO?Y�E�����rp��Z�t1�m�6������3>1�XQ�-QQV��%u�_�9;x�l�����
%/O����>ew[�&XgP�B���"�$hS�	5��v~ԩ74�<����Y(6{#>�	'�.���VD킳X��o:Q����0��ܙ�-#
NɆ�	ȃD��H���;��zs�@�|���o�Fg��'�Eu~��(;��?[�u-%�\./��Q������r�k�϶t���<��ݲ�d�Ո�57�<����[��5i���Vb�<`Wj��tj<���d�Ԃǫp��1 ��m@�uQ��� ���IR8X���T]�C�ÙEK��t;�g��d>ա"�����-�7ݰ�<K�c+�!��Lq����y�}���D��B�����<}�<�;�K����L,߰��G�Br��JZ�]	p�"� �t�u}�kw��+l�O�R n�ų
�u�~�a����y밠q>��a�@���=p�t�
��G�C�x'w�·w�L��<�d#3���j+�۲#�DŴ�`+�#�g5�1�����}�{T}J�)��@@Z8yO2�7�`�Ra�����=�i����U� o4�Fq��Tզ�:Yvؔ:��,��X��|G>�4s��BK���Axs%B�"�h�O��L�<�=�Y��@��ݫ��:����s�	6YK����$/bp��n�;�U��p��kA-B�B���t,�.��u¹o���w��;�(	�9��Q�6xe�L.%���~k�WK,���܋�H͊
`p���R g#�Bπ�½)Z��'A��P�Q�d�k���p_q�Hp�9dc��mD
je�52���_�?��KZē
�%�j$�1�D�!�����d����w���)����jT��������
ϼa�@���~��Y
_��*�l?�8��bV��\U�$D���o*�-�@�W3ֈ�v�ߑ4&�<c]�d�z���K�Q��YQ�e����GtN�U�&�28{6)�ƕ�O���y_�yd��S?�y�!���������^�%�7����z�(���6����o]/��[t|�@K]T�����G���)\ǥJ���(�I&���bZ,�Y����RO�_6�L��ۼ6��\���zH�	�~�]j��E��[�6w�	r�a|n<�2���4���E�9GΪ ��Z?�d�aN����]��{v,P�.��%�L^{c��� ���ԽϞ��o}f����d�d={���5�mM3k�N�0�������p��~��w_;�?S�␵��z�D��̫	��ŉ�cw�n�aVzd:�4�o��ñ�[]�t9�}9�Gw#=�������Ի"��3⃱
�C��V7ȯt�L�Oi����p�9�v��b}e�\���e��+�n�ɓ�.��p]�]�Z�}��~��P:�A.Ф�ZTsz4�D��3ġ��ps�e+x�z��x7c���3vS�q7�l��Qb�%G�U�C.��X����y�^�>#�?[Z�]��_
#"���#s�����;2����?땯����C����㍽�#VO��'ⲝ��>�Gw7�n�E���%e�de*i��A�cc��v��X�ϖg߉+cH��D�A�G��p���)O�J�6��]�#���"&V�Z�zԕ�����O�������l����]��7�
�M����d�|�a��I+��K�I��x�*���nY2�آ[9�J��2Z����{��@�sl�㧉�p�N�yN�����qU�{z=ru����8���Ԩ<"�����^��w^�Y�'f�*����9��ml�5�X�Uھ	�|�T�ž�l���`���e"�X�3��ن%��	���d��a�.�Ņf�H��)�ʥ)���$��	n��ݷj^BS�d�h:��Ъ\J�e~��3�i��q��?p�s�-ꊣ�BD�Ȧ��46�����:���H[�u�h�ǖ6���Sύ�Dʥ¤�kMfE|؍a��ϔ���"��u�� |��1h\���ii!s��7X<���;�vޤf�S�d�dy����͝<�����uŨT��\'q�3��hTIUt����5�)���z4��`r\�:i�G����v�����fD��cTp �~H�����m~*h���6&�
�����>]�����ŌG#�Y_��^D�D��[>���z��M��)��������ۛ5i*�太1��N���R�d�����?<��4�hI��7{�G���j�= $����r���K�n�(3Q�
��6�$��՟z99+l�w��~y��q�wCu���ĉ4��3�_�o�J�-�$�e�r��aÛ^,����"*��B�԰�T������'�]o�EFK͜���E���c�Þ��?;B�H'u��&�X���Mb�;��2�B<:Nȭ�:Ǧ�tέ��>��is���J��ê�Ņ�����T�sm~�J\���Me4��׵+�֭��D�N���EI1��|=m]�9U�1!F<����Vr�C�(y���]�jG�o�!?�k:��Ξ�?���p�l&<S���m[���ň-��=�K(l���İ}�7��#O~~Ĕz��>6�̽����(`�i�q5�~�>bW���fM���W��S6]ɺ�� !	�.��s���
�)�X�Y�D����,��EP��X�i:�b���H����w6HV�p*��O��M�T���5#�_^K�??J�X,����>����Ys�n�����o�i#E��.Ok;TJ��A=es�G�a�x���I��!�P%���&ɰ]��o�%{�� ���C&5���P�V>���j�c
)^�H)�N��P�0U�G?�oX(Y1,4���6ʌ�S��k?��HkMs�T-����p����C/�QNb,�a��kI��8������B��9�]q����HB"b�K���$y���kkvVrbC�%�[�����6�ȑN1<�i !L��`J�"s|��,YI2�T�FK;K�k�<I�ї�q
��̄��r7�{������%�����<��mc*7c�i�l�i=P:.2����l�fě��1��Ǡk���}�6O\�L�D�O8<�Κ�U/-��zy��P�|��mNC�|�
[��,cp+{�b�����~v�������!e!��;� �-��j��޽�<LO��ӍuY���f"Ya�9��Y
ᅹ�"��:-����\	�����s�����fN�����d��܌{�����5R��}�k���=�tm�c�+����<4	�����"S>x2���/�!(���rR���Pn�����������4���X��9t���6�7�����3�Ju��LT���觊���$鋊+6�	��N5�k�+��[���EsdhK;���]nˇ�<��ڟ�y��6�ii��R���_>���	N%7��uԅWrEz�gE��&�U���-l�)o	~f�2�%��*i�#�rB�.x+�����`KO�<��F�q��ܛ�uzW1�T߿��s��͟���u�Uhm��c�X��#t��jbz��ۇ4��~����8�r/���-���/t~<9zJ�a�$��TW��w,�Uͫq�{��綺��}��V��6�OX�]�Jp��*��g��9�XD�`�������<�iU:܈�6O#l;�*N�w��+�' ǽ�㬙~T� �l*I�\�NyBX˹!&8ޣ���g��J^9���~�b��Կ%غ1� �:�V#_!��X�����<s�0Wlľ5� �
|��2h��~1瓙�xK�N�����}�F=m��_w��˷v�D��*� F�a;��& ��o�nL2D������Zc�T���{k7_�a�����h�)̼����d�R����o�sC����Q�2��r��I%=I݋E�u�H�����8��N�='�W5�s,|����Ì�	�og�y�H���%?�M80`���e��I+������1�:R{ޟhLj|�=��Zd{mz�����Y��PS��I4����l��.)��U����(5y�$ܤo'�챫�^>���X�z��X𻶕��o�o���/���O��9���n�l-�9q{^�]s\��c4�U�ly�g�t=����:5� {	a�sI���̄roZ�{��0��OjP�9���j�Gf$��ճ��y��~z�o�o}I�� ���6�-��&&��:o��eU����z�_O� �}q�L���󭟟?���?����?t�1�,lՇ��p�i����{J8K��ne�<\gx�,��d=��lv>.��l6G�R���3�u��JVI��c���r�K�(vqz��/�;��ۋ�Z�&� ܏t���Ǳ��)
�?>fa�����\s0��E{~�A������\5��[��#Y�d���Ƌ�Ze h*GZ��2�]*c@����?g$.K$�j��o�b���#�kt��[[��d"���2�	�2�߸�أ��閴ħ$+��3��-��ع�+�%-��[�X�X�薇�vˮ�Qy�ɣj��ҩ��ӣ\��Ģ�������|
�q���z�D�Wa_
C���a�2�K�Ƭ8�;K-�z�^��Yv��K��rh�� \H�A��"�oӺ��/{yv#>�v��Jf[�Ī�
��Ӏ�Usz��v�wO������>V�T����+Qu�}�c>�ݚ�f,�|V(z��� �\�=���B��ͼ'ѻP�������]~r�����B0��_��	ɤY�Z߷- @a\#��b̛�`��ug;�#�e����K6P�XZ$�=gl�9�Wy�Zu?��,;U�A�-���5���F�+/��Ǩ�����f&��L&�3�F'��7�!p>@:8.��/\���
A�'zW Z:,o�>=�>_�p;�?Tר��熱'�n�Νk���b���%R�c�m)X{��1�;W��g�`����7{8�4H93��>"&�u�p{�������H���N>��}JԶ7}|(L�L0�F&b�ѤU��M����2������W����N�y4���t�}dB�3q�g^�[�؆]��:��Δ��尻������N��1t�%�q?�a���-�60Pl��-���)����asĬ����b��m{K��x�]���(k�%���qF�NC∼���C.\��$)/�ޓ#&��~6��22
֗ �l�e2[����ȂO]s�hٔ?�,^t�`>��L�0�^N���\�~>�c���I����EX��t���g�~sl�,�m/᭽��p�!��F�G����!� (f-\Ź	��*������f�)nZ���C�Yg�`�+j��9C����;���� ��a(c�PҴG�3��ʁ3��m��e���@������t�X�Pg��%5���%����Ń�~��%��  ��@�\��/����3"~t��EBu�49����E5֬�4���v]��&��z�\�T Yr�{��g=Ք5�}�\������#/��qd��N1>��6�q7׳�p#6B$��oeU���R�71	�4�]�,���j:'H�{Crh=��P�Y�.V� ��l��|LI�%OJ����5�eq���w;��$�y+�-�r�z�zλ���:�`�q�U5ԩ)�Z�o�)W@���u�GKP�t9�z�HA��E,W�0}�WO)�}G�hk����ʫ��6�K�ݚ�3[+�ȩ�o��j�J�)eS�M;SF��p�l[{��{,B�ƪ���'_g���
�+�	@��|�:��ݧ�K��+7�S�hn}Bp=���o�.܁���> �hH�����;�ӛ�r�n�jL����[:��b�w_�;Y���+�,Z��\Z](�,�×��DBp6�쟵�w�Ѭ��8�ys�ק�g��T;���?w���q���2^AP޹_$��"�W�3�4���M���{��{G�&RlP�����F���r_|�=�`	8����wVP���������40�K�}}QGl��-�<B���'���/	@=T�S�l����	�sy��l {�f:ro��X]f
�|����^ңJD���OZ���Mg�� �_g "Q��CPg{8a��z2d�B�?�v}�K�a2�7�4����?�A�U bYf#���痲�	��N�g_0�X���Iߏ:%�w�It���3|�/���o�(q����p"|؛]ƿ=���@m����;��-ա[S���yo��1�S���yNJʠ���B^���W�i��Wf.X ϩJ��hcQ9�ґ<��m5�J�#��T��ݛ��!��
�&@:Z%���+�BK��K6����l(�X��u�(ݝ������7b�ջ�P�g��Ͽ�x�@���c�䓴��?�o?G@¥��e��O6��#������U�Y��C�Xo�el���'t��Otiqa.���)8J_��l�#/v뺃�����g+c���g+���5�G*02�6��c�E�����)��Ap�5;�����ؔ��H��o�����Y&�=1��m�F���M�}�=G#��`b����׽�ϐ��q����2	q���v_�_��(��O���At�C�/��C2��W�k
�i�|/[6)�gf�:�z�;I�&�!��#��?b�/�������V��O�a( +��<*�ߠ�rz���9}w�e���m����k!���kYc띈�u���&~8�3]����g<y[ZQ���~�e�?!�o�p=�{JE���b>G4C��Mc��/��l��G�yR��#f�,%�����g"�Ďy�� 5�i��N��[k��W��#*��kNr�b���۩t]Zz���ݳ�
�V)���Wo�L��zK'�n�>��	��_k����%]8�E<�Xo��8+7D��n����jB�\V�'rRԖ��ZPԨag=gE���;cq���~6Y*�p��1�U���nބqM��+wZ�NC�j���HO�m�� Fz��]:4�a4����묇�5��dM�0R�W�1]b�4�T��v��:��r�k��z�T�Cu}S��h����VOyT̔��8�! J�ƽ�Bދ��I�:s��y;
"&���WiԳ|8v��-��[�!T�I${6^'��Q���[L�^�v��,7��|������S��F�&���2hO�U&m�6��@��Ĳ��AjT���A��j}��i��OP�|]g5=Z�}�^����:a��������{f���)� ��x����7]�a7Cj/���s�`Ȝ��'��%(�n{`�ˀiw}#Y�#񤄃�bS��J��]�f�2��a�u�Э��c5���\0r60&�?��{�?s�g��5Z���P2���4*���)x��j�z�WW(;}�mK�H>S;�dwd�q�4�rr���M��႟|cG�酉չwx��1e-������E� ��6��`���F_�x��g��]����o�GR�4e0�k���o}x���W{5�;��C�GF�:n���/�'���Rl�������j���r��a��`C)�B�/E�'~�G� ����Xi �湕���I�ܾ+�&�T�a�����@��>����e�����8����xz�Xz�Du��Fvl6�tY�J5(���_��RȰ�4ܪOp�S!�:r��M��ũ�5�H�n������v��2���.OuH����xn����Q�ϙ��w$E"�y�J���_EyU���Y��UDӎ�ED�;D	��ԍ�#�2����r�Djv�y��DOk��s��}(.vG�g��dP{��W�0�=�c�>��}v�C�a	i�+�uqp:j2M;�zɗ�&���J��,�)d�x����l�X�j�8ůn�����t|+��gSp𩘉Hw���M�a[�^���i��Pz�/ه�S�'�\s?k��N�#�3���٬qO�-��iӃ_��0f�B�]g��_����ʨO�����b.Y܎��
����A�pT`�qo�Ri�1b�����J��b�i�®MF�H������)6"�H�!�5*B$C�2zI	�#�|*q�LJ��4��~Z�O�2��qk���cj�8M3G�ӌ�����eg+��~:� K�X2筝M��bI\�QP�u�H�����LÌ���}�kxp��*���^�3����g�4w���w2�_��N���ḇ�	��Up$|�s�����bHBrm�����$2.c_@��򞣎4�~-���\ќ5i��w͗jPGTQ�0Fpd��)A����[#��g�.U�_8Bߛ(Eg���־��ģ�����LM�v�
pK�� �}i��Y#*���v�u��?�Y76t��̠g�R���{"KŨ�'�S���q��	����~/y��">M�`��F��,I��J�)y��Z i���k�wo`pl�,�vj���\�^9��#8T�����k�����(�3�r�V��N��<�`����#Z��ŅR]1�.�,@
���7�/�Q���"�	��Vv�L3sVQ毖s�r�o��w;��Fe������\�zj�(�VY���<�"zS�n��C��݋����!�+X�>��UU8(�^af*��%���M<��ޑY��0�.��jMW�)�=���c\�b]�f>g�1���+��>�<1�K�*�D���C����sO>k1(�w�M�E���$���-�r��f�Y���<�F�m�=�����	N.��u�J��c]�8�.�K��Xg����-_��&J_��SKS��*���Wv2�뫰?��1u�M�)\���Է]1"U6q�����(�sZC-�*礂п���g��/T�^{ƞ<��UË�f����?�"ס\���*�����eU��`�ΨBZ�����O	����;M�w��4�����!��o���çYQ�(�hǢ����?�a/��~�j�ߵ����j������cc�&�ʧF{R݄�{��b�mb	^C��Jխ�V��q�AUp;Gέ�^K3�(ݭ�z.�#����y���Pml��<y��Q�=���+z���MW}��Z��#���p�(ԯ���U�*"$��)�"�ԃo���O��Z����ݡ����~�M:dY9sȯ���2a_91K�!>��Z�s�q!��q7��Q�z�P��h����~O�DbWt�vX��K����/�}?|%���I!�ؽ��}�C����M?��!)T�0j{oRR�2>��N���Q�2��I������v��N/&T�)�GL�5�j���X�iA.�Y�)�Z��_i�7�"S+�U{�V;la��ޮ�c�3Bஂ�l��MOk�FA�e})�URC���1I�ۂ�q�OR�V�\/'���%��|��v��`��\E�V����	��Wm�*�i���v5�ef�Q�koC��j��h�_DF�cޖ�����+���S��)An#K��*�R�jiSF'�[�;�}6���³���9Xr��'wI�W���6dE^u-7IwH�k_�o��[+�D�n�c@��t����\TUr��e��_�ԓ3hF������w��	�ղ�h�45V7�I<"�]O�6vg�VP���_T�Yo�j{;i�)��AO�=��*�nE�t6Q�}�ۛ��q��$$�ZE���1��}ٗ�=-g��d׎PF����VNR���dO�Q���`6�(4���6�U C=��	����7�q[�E�-���=k;
/�4�nf�8Xd=���̬^�xW�iT��֦{�]R&L>�lUR(L�VS��Цk	 .���l�A�ʳ���>M��6�#�z��R�p�,�bE� �Iҵ���=�r<��I7D-T��s��X>z�MG�>j�j�O�+!W�0��5��.̝s�S��w�XG�Msp���ȝ̮3�k��j5ڽ/3��,N{�����7�ʏi��W�I�5�7s�:ǧ����=�|敏�,��]��L��~�S��;�h*�%�=�-K�"Yvh����ʿ�~�}ӥwh��޻�����_��S;�s���(�.$��w�854��Q�C����k���f���V6M��]���$�g�+��8xL�NFN����;�R1�4��=�Q_������=:<H�%��~�v�������x�c��Pݣă���hni]�|����+��=�|��BcJ�~����a~�5آ�4%R��2ZK�����R^[][�#��=�FE�������{���	�*�����_�Iy�׭�6��%�A\�Le)/a�9��)�/{w����%oR�)�	v�=�d�w���g:��Qj"@��:�O������D�UI��id�`��Xn���u e��@�����W�Wx�+�*�/@����g�B��Q7��7�y�W`ޓdƱ����c3;��蕘:� B�I{��~�~��޻�`��������X��l��˫�>x�Ζ�(\:�V�Se��pN��V��v���Uo���\�.^�yO�Ց��>-]M�$]�7zq&B��YK� W,��-��EmT�1�k������A���Z�88o�I.y�CxU�W0�5����z\k�|��.T��${�L��fC�r�� knQ�'T�5~����9TC��p� 6��.l,{�c� n�?���O��Y�E$�Y[��CA�J���%<�u�5�H+�>�����9,����7�Mޤ�z���f�����e�:�5��J8O|����2�=��kU� |6��j�XË��adn�~�����M�(�a���Pg��C���<D�� ����_J�U,�i�����f9<�5v+!�D���8������zV�[�k?�>�<S3�#��c;է�7��'�Z6C��$��u��M'I����(W]I�p�j�3%��R7웣d� ��_`�Li��|�6�sȶu� -�v��=��o��s�����˽h4�����_��j��t�!o\g��b�c_=�ö�D����}���9&9!P �Q�D���w���(�L+��׺�'�k�0�`��Z��8��(2�zB\©�2��)��Ga/K~;=���c� �A��~kdl�TT��kn@x���y���6I>8���)B��%3F�L�~���xAK�u�i��N�H�N�<��;�@5��~�q��?%�EX��0���ÿ�[�^����w/�D��`���J�Oz�����(����p��X��+�ȴ�toG�rT�6�%^�[R���?��oL�qe�rO��n�d#�7�K
�0�V���=�߱�	������q�KS��������0�-�tk����E ���+��&ʙd����ߓ�R� $f�ץn98�v�~+%q@,���U
d'���6�Y�����qw[B��%�+q�$��)�e���o�E0�c[���ń��R~-�5��*}k;�!v;j��ߋ#��D��3N��2�o/V?�V���8���0>��;�C{�."�6i<z�o_�MF��
&�0?e�u�&Z:{�e$�5g�K���S����Ie��O�Ͻ�<JZ4ISc-t� h�ROK�)�����M�K{*��yQEPH�K��d���s��i����g�x�&���k���r 7)1D�	1-ܤr�����N��}@�mQ��܄2R��ڻ��&�\o}�ߡ"Sk��z*c��w:�Q���=�ǵ��rV��#�D��B��ᕢ��f���ұ����Ϥ{��Tc�cYM��E{���x>??��5~�k��I|ff?��9����$�b�=�#!@,xzǖ&�*B/��V�������'Q��'=Q?{?�~����������h-{8ԩ����q�����q�K��un�斡���ESW���nC� ��{�f)�j-�� I�c
<���\�˵� l:�{95.��C���FD���:#μ�ߋ�G@H�ղ���'I{9{�PS��L ���K� �	P�:b�ݏ���(R����|si�K3~�յ�}`�zK_0�F�+�:�ޣ��b�R~-��މa��p��n��ޜ���V��aZ�����.��X��ҫV�����F3š|���%]�L�~E���B �֪Svg](��7F�ș4x�!y�~���� �KR��eﾯ$�=�#���e��Xk	s�R����� I�Ȱ�W���Q�§��Ԩ��� �(ة�����A`��t�o� ,+��-���E��$���ޫµm��m��ȼ����J��g����Qu�6VMR�����dH-���փ�������p(=o����~},7�_��`�7#���Dzr�ױ�����Jt��:3����M�UVdO��U��H���+}{H��g�]])��:�o5yW��n�Z���
~?�3���h�@���GX�յ�X|�_ą��M���k.�;�L��<�4����/�d�x+|�G9p�����LNu��%J����-U�
������ab�ELQ$^��G�	-�E����U.[����ɛ����(D���B�i�ߊż*Q��*x���RzA>����b�C~�u�y�f��?��>S���m�s/4+L�D�qRU��3�������ϬQ���e1/�E���	|Ƴ8��*<���~D/w���eumY��щ��ٷ�b����]k��͙�I�tnm�b�]����3�u��jjJ��P�хG���,{�ܛ5k���St����-Q�����%�kH�w�O;��!Y�be$�5w�ܷ^,>���ˈ5����un��O���.���b��}wc���N	�h}�[%��\4�����2v�La�U���lU��ն�^�G�O9,l�c����轹A�aN����B���f�I���6����1���������.'�3�L�ug��b��ř��6���*+��k�#�`�N���T������0�Ϟ�ƟJ���3}�����������L���PL����}�g<�	]�muϝ�Z��w>���ot׿�G ���?������ ���7ٱ��4���%$��8q��_z���;�c�w�?��{T֥�z�v)/Us�֍}H%��o�l��x�Ԯ��d���b���d�L�O�gB�Q���2���G���ņ^ʁ�o-�U
�����3��J�S�LQ��e�?w�gk��&���[z���o���� �f:X�$hy]�q�ӗ�g	�0�wFT�+�3;H�S���G��$����Q�w�"�б��Sj�3�NM�׍��n�&W6U,��U֨3�(����%���#�ǒzo/���Q����mp(z�+K�:�ܟ98�_Ӭo%3S���� *�R��V'&~mə�[�)L�1A���8+\��NY�.�9,RK�n{�v_���~��:�b�_`l<`ȤcP�b�dFUH��X��!/3Hf�v:l�p�=u�l����3��z�J�����Kvm��#���rgNe�މ�0�-oa�����#&����;�1�=CiZg�7-Gȓ����%w�����o��L�i�FP"O�Δkb�R>l&Etx�#�¹x0s���	r
_��X�M�S�~�U�G��zˆla������͔�)���IeD�\ pϛ���ޖ�����ΰ��H��g���ي�s]^���r���Kͱ�7��3��շ;9iZ���:<�]O�Ɂ��axY�5)r��ST����a�kh��.�,�u!<�D�d
��J]D��A��ڻ@魳��!E��7�%V'�l�_�{��������+>S���������i����c�8C'w�\�����/_x9R�⍌��n�xX����]��-���2v��� k�$��ML|�Lrxa�;?<`��j��?�2ÞƎ�hx���U����ͼ{��iM�ᑼ��P����
P-�.<�uBz+w��9���8~�۟��<�Sl0��Q�eB�7;��wT�Y�7�<<#*
VP��*EZ(:"�Q:���L�Pt��JQ� ��HB�t�AZBI�=$� $���� ��q�Y�;k�X�{_e_�w]���ݱaj�Q��%�'Iu���wi0b��a�+E�b��ĝ�_8/)3��7�h�Q�����Ѷ$�����sgGdz�0:���h�l��ώ�ZhM������f^���|�NQy�h����e�+�(�_��f�lV��[5/�������풬�nN�,�����ð;o��Qr�.��4�4��iΠzZ$i4���h�][u�'	�|[�j�ө�9:��Y�]NMu=����������P�;�D>��Zw]���?�z��m|Зc��*��v�����D�巍@�x���D�)ԩW����z��AS��H��d6`�q�F�x�5 ;͊l_��(Y�|=weԦ&KK�qY�����`����Y1����Ip���<�@�W>��N�D��>�,��3�o�+P�u���/��.�]ȥ44�}�Z���H&b��z+�m.�����L�Hw���v4��<9+�W�d�*E� �2�������]v�mE�F���Z{[�K�s<�� �K�n��|5�n����@Qo��-���f�U7�[rJ�Ԩ���$L��8}G1OqHFf��:-.Q^ѓ��?�?�"��,X$3�d��u덖��l��a����bn0�`lt��0��lx�:����������CX�x�&d��E����RH��%�!N�S8ʧ,%�j��x:$�:;�
���;{̬��ŧ�.��~����z'G��Z�W3�[C���Ӄ�^��l�|dظ��ʒ/D\�y4x��S����UO�g�J1@��j�9Z��2/>-��v�����%p�&��7H�#tRWɜݮ�;�K��T���gb�c7��������\���ni��Upi���^�
+Z��x�.�1�q��g9���ۄb��/�aĖ���2�WK�T��5����¦W�'@�qY�7��{����b�m�Đ�:��dY#���x!)he��瞇�e�g��0*G5T������:eF�+��Έx��.�;��7�<�f��*�Y�lwp��zZ��'�e0̊Y��Hv+�#��j5�������^���j�ZW�-]�$U�Zy$r�п���
Ez?c2�
^Jq%wr��=�Y���vr2�Ś� �ז�1��	s'h�-�͞����Ə	�s�4��V"'��p���/%������?�;��U��7��}�����]=��ld���C=�f�Kq���GZ��������;*�F�i��O�B����$ӡ�����!/��6����,�&���Е�>��&��o���\4Oa�9H�t',��77�,�~��]�rX�_bI�G	��X�4�(�e�����ӂ�6�Q�E#n�P/�>{ďt���M�w�~�E��:�l�t5��(։ڌV�ռ���{�z��-X�y1*7����?�oc�|��R�O���&_L��T�D4{&{'�\��;�T�R⺳�`���&�Q�6L̲ƶ.�b0%��-�İo��4�0h5����)�^>v�H�W��d،�Y����E�c�m�-�����.L������}rr�{(a�:\�Nq᷹8,G' �dbK����]��vw�j$�03-�8�m�N�Li)?�HQauvS��͓�<6�y���|�P���T��{��iC'@��_[Brs\,A�kbs��C�Rb�i� I��t|������LF���X�5�.܌ 9,��V�������nC;���7{�x�������(V�[n���|Bh������j��u��j�3K�ylol>�����kc5q�x���]yzS����n�ֱ�V�%��}+/V�� w�A����R=�8$Af�����t�,65[[fk�BR�̒��FPgQ�Eu� ���u	���(1w���-�c����¶��Q���o�%��i�-��I׌�!8��6��B��k�N?�����%i�jʒ�����%�'��6�'h5�Eɤ{��x&a��ȳ�Oh$狡Xu���;�J-�[�3�N�>��g"��	@��Q�K��c�m�6^"�1N����JR�&רȟ�T�pO̽P�A=�"
��k��2���w�0~O"j�{�A��9K{b�p�I�a�*��
�އLH���A\6~������6�N���.�T�b�B���JN�>/0�;W��8ӳ��v�i9�������7�0���r��;}ۡ����E��w���Kd�6���o��Ռ!��6���뽝A� 4�,�ɘ*�,��BP���cF�ي%�ʋ$^��<�E-
�Z�R�;Cm�R�c���
�p?���ufaH>���l;Xg��6y%_˄�׏x��A�Գ��JFZ��/�2�Ԅ�̓�b��'�5쨃�5;�LUh�3סg�#�H��ck�H�b��B�Q&bT]��NŹ�MX��V<KI%�%�o��4db��D<iݯydk�(P>�LnKY��;!"��4X6l�v9��	���G�A;����:�`�-6Ll|��;.1����oE!�yc�����=8��q��]���cA�ٻ���BK\Ѐ"�����n`h��V��	��S��\�9�*F�%-ĵ�.z[��N2Sy5���z�4(8�v�'�%R��_�N"��ǒE����5�	t�U�1!8�I��D?�~���NPLg�nyw�:�wڰ΋jB ]��R�aНB�`�q����F�I�aH(���|@դ!���5m%B1ld��Ψ��5�<9��<��lJ�]m&�m�6�3�^:{���P7��vʲNgؑ�eW���̳.����눌V9͍%jtT�+;#+�FԐ��yq��2�"z{<�,��e/��¸.�CIC����R��ؑ:( �W�F�p"��������B��"-�{�nkh��y��Zw��i|�v�PT]Y�� (�ejaC0{�qW,��zAX�k*��<�I_����֯uf��"i�&��S���0�;9v&�t�n��^�z��u��ۉ0�0FO��7W�s��#�.�u�"-fu��Go�
�2B����� Sˬ�5�u�����H��C����؛F�C8�ۡ��Ob�]�Z��)��R���803��������	���_��Nz�"m&����y���}65��*6���{�3�F�u�QØz�н~Qϯ��>��`�(����E)h^�����e0n�G�p�����i�&�lB9h+��;�έH����=������Hܛ˫�y�t|H1Nq�rWF�u��	��nL�r*+5�VG���,d�C��/�yb:[�x�1�r� A`���2x�{r���xs&CP.A�� n����a$��+�˦�N�JOp,*ǹ�,i�!�B���\���������V-�gp�PȌXߔ���I���`ހ�г�XB=3�Q�r>�a�h;jŸD�U������	�|�p%�$o h�+m�/vapS_�\:
��Q[�p	�e���6�x��4�1t�K@[��%@�L��n��@K"z&�+�i���/�=�mM���yxs4+C�-�]F��&D�z`�W���Έv�A��mt
1G���/�.�=\J��h�j5(��b���j`���}_K��]ص�Z5/W|���$q�:�
�`����m��V��Wc#�D�cZ��-��x.�ʩR��}��'%���l,���`g׎��������U���
�����?P̿H[�������ߔ�Z�~�5�P��e�k�I^�]z������I�v���Aʿ��~f���	R�v&wX�?�6)*X�&O����^\�&�{�����v�� ��B*���/C��?p�M��z"�	����q!�*X�猨p��R�[GX��Ϡ�s�6rz�ˀ�����bq�9�^p��ZeHF廵ۛ=p��;�v0��@�ءt����WŢ�>�n*�)����w^�����ڀ��M��u���2H<KXы�\��ݨ~:��P�6��ɄJC98�,�v��':�#�*��\A �(g���b��<�ٶ�ȧ+SCdM���s�)�x�Lb?V]EmL��>�|)�Lc���a<��2��
L�Q<���5~%�}�O��(�P?�������Y�:ٵ�6����@�}�Q�׆lf�K��u���EKRX�eJ5���0//ϭ�S���	-��	G�\H1�=�8h�c�5��U`��ow�E�j��,_k��'=�.|m�\���}Տ��g5�|�1,I�g[ɮC�Ê	wc����Z���J�&�6��i���RB��	�mm��|�Vf��kN�m@E5�ƞK�8H��Ϊ?+MTh�R��#��z�r��b�Ü.����WY��d�N㢂+��,M��DQ��>�vMsЦ�{����#>�u��?�WY�㘨G^"-�m���]+�ou7���S.O<�]�6�M%�BW�� \�k.�C9���������h�4�����r�E���ej#�#	��H�w6���V��/��!�� ���~�l����4?ҏ~�� ��LN��pB�m�QI�s9���b4`�^��E� ����n3�/_���k�R�r��zzg}�#m�,�!������'%B�����HB�� 2�h�M���8w��L�h��A#D�(���Cq�}c�w������&Bqy�����yx_9�w�������G��d�G=�.g�D���f�z�͕��fV��.�>*��w���\�>S>|)`z~��~&�7��L-a�]�����z+�C=g�����C�Y_��b��&��#�Ҏ�^���ŹŶz>���w���
�aה䩁[��u|(������-��鵅[�z0C��gk���<�F���I2�p����~���Ca'�;xxd�7]��1�ꗂ(ȿ^�}�[jw���9Д���"�;�<Z��q�k�k�B1�x0��1���l��4`�PC�����QF�o����=S���M�~�1B��d��C�)]��S[=�A��#� �_F�G�7��{��-�x�YU��X�<����#{d�'W?�Yu���a���{Wp���{���V��:��ьwR,e �$��mD���.t�}{K�(��?ź=,����s�� ����Ә��HO�KG�W��=>?:�y���x�g�Yw�h�T�~]GІg��������&�c�ѕ-6~T�x�q�U12z!����q����4������<�ժ����Q��o)����Z�ܷ�"�%��+�i���������e_U���>6f�W_֥�N���Q��.ķ+�wng��%Bm_����2�Ym�u��8�-3��kM�~��(�D�}�O�!�}t�孝�Z���)�c _��6��W���>j�.�S�Dj'�|���'}Ի��<��$��q��
�9Ӫ�1z�!L,Օ�����]��V���H ��E�ћw��{��Lz��(<ůORZO��O��)���w���+�8���$oس����U+
�r�^�S�D7�s�Y8�u��������wT��r#�Mk���*2�0��9�ڋ���un���P�T��P��o�z�������MM��{�(��~�����H�G�dɱ,׸���}�ȱ�b�*d��I���]��;�^@D��vO���~pujN1��]�B_5^��4�q�OYI-�~��k �!��I�U:e�v�ƒ��Q�\�>��w�]� ������9�Ԯ�`g�r䥳=
A	�M����gg�_p��r��O&x�9�X��g2"lz�mX��So�<
Q/Ʀ|2�dj���"І�E'���C~���+�	V�WPL#W)U�3Z���A~ rKʛ��Ƣ�PS�.KZ����C��[�f� �p$��I�ZF [��w�([����6�,P���WF2Y�� p�vQ�o_Z�nd/u�NR�¸�I�B�i�E-������)Z5���ɐ�������{���'�h�L4��/�"�y>ҷt�n���#����ƺN�Z��C~)2�m�^��6�OPڑm�� �%�|�\(��� X�n+��;z��Ф���ԟ��5�]�ҡ�Α5Ė~�p�k5F�s���w�o�)IV��W�C�]�g�-!@�)Ԍ�{�pۦ&`l�5.�.>4y/M�w衅\uNq��$�e���.{�? �����TQ����w�b��8�9yJ�/��#J���!�~��=�~9���(j��7וjd�!7t�h���&����Z��  �t��:-�sKj&?A�MS9:J���?7�`n�K�o��D'�`>�ԟ� 8/�.����E`����_�&7�0���h5������g��:�@�N:�n3��|�qz��BG� �����00;_�bJ�kq�åC�`%�l@�2ؙ�3�g���Qנ�n?%Y &e� L�Ia�t]�mfc�%�@��^K��- l91&��/����3�7]�4T��jK�z(�z }�t���t� e�<�+��M]�b^��,�)m�[x��>1D�Y�v���:(����m#Ȋt��ZY ୤���~'�,�c`�(*'u��k�ͤP�{Z�����2�[����(���G��٤H��x]L�(C)���^}-�s�̯3O�,v1���{�/>��%�k<�1T�U��X)[�,�.G T��N�P��,��Mho�����+D��W��XfD<���e�۰��y�`'R�K�	6��(��0p\0�����{  ��5}a�伝�!c77�v?X�V�}C@�XHt1��s]H��0���v�=�V��t2@x�^�:T45�W�Z!^�U��a2���
�?}St I����.1Ǧ�e����e����놀�f�ѥ���}�ȗZc���jZ 	�x,\	��=4�B��؄�~G ��;M ��0���LM��Q~�X��`a�m�y�hf����wޚU�r�̃H͔�$�k>�3ʳ��4��i����ʀÊ�E����)�[�gk w�'-J�>'������g��t?`o^r֎O��(V�ō��  �9m�[,���C�	$r�t;��k� ��9#[�z��Brl�M�1��j5���н���w9L*aV�Y]���E������KU>��h}�vwW�􎇺k&3&{j��.�W�И�͗���ǔ5!]_S&����&��hjG#��^��I�ۅy�Z�G��;^tKJ��P4@͡ڼ5�KR�	 F7�=��	�7W�L�>�la4�~����B3�eg������z�{屋*P�����^0�♸9ͪQ"��չ;_��)�D�Q�����K� h�' D΅"�d�G��� ������ő���'9��p��Y;M�e��P�IQN~A0֕����s"E�ʅ(�.^P�= <�F��.a�|�y�*6lcN/�˲�,~}X�Z��r�M�y�hgi�;@�g��w'n�����B��^��F�=�0K���;�-�PMe�yT�*)����pfV���maDanc���҄�6���+4�e��KGw̱�3Tp��kO
c����
t�M�]��ʴ��	�
d�/��x������m
Ta~c8mJnO{��η��v,nSY*�I�%ۖ�,F�q^,��~w���QM�~�K�
�T���T�@� �P�d,w VX�l0�x.|��a��P��22[�35��K���/��4S��xA�r���vyC�2<��X��"zV�zp��q7���}�#�Y·�?�i&���\���`4�]v;�E�	��̕"A�'Fc�vr��q3n`Xq�Z���(����⧆/O�_����]�������wsbH�vO���u��B������	du%�l�kh6'Y����V��-u��$�`�7��Xo�"A[Xi��d�o ��t_7΋F2>�A���6, c�r�hfE��fv{5M�c��Z�G���	���Rx��Ii����9�hjl����/���k̼Ak$Ԍ�L\�À�IN�L�Pm�xN��r�E��ȣ�F�_�!��w��$�B,3���̛�	U���Τ��U2��f�:W�!��n���P�+�(���������n�k"�� r�e�ʂ���EدXK�N+Kt\ߞ�n��Ҹ���v9�a'��3c&:�*�6�3�=պ�赭�fZy&����@	�:���jlP��������-�>�W�@x$�$�]{P�ڍ���QY��0}R�-�VH�����~Ҟ��W��YE�&�8�8ɹ�I�AS��&2�b��,Pj�<��O��dT)�u�-�w�,�[nJ�� �n�T$��/���c�P�Q>�<��ϯ���.h� 1tM��2�d��w@��5�k�8��h�Ch�jO;_����㺙�/��/;�&�V���>ˍ�W��K���w+�s�f������i��A���!%	�}S{]�o*bL}#+�sVΗ�Rc�W&��N
�7\y1*��K���Z�}=�^�#�M�Y����A1�}ۜ�T;�1�{�����\��<�#�^�x@�0���tK���sCA8����Ws�o|K�6xj�M��@�cKoל���IG|>����1�}�C�KlTKʡe�%S���$g�@m@�H����zLA�d,�|�>�Z�ԁdyA��1Kd�@�Z�R+y�l�	O���?�;�f�ܿ�T�s7#�CJ���A��*��9H���"�����s�����ԡ�(z4��&�y/��|N��<����n�/xd��9�F`�Mѥ@��(���x�0���:(7Gӷ��>��^����\~�Q��碛v��V�΂9���Ea���lR�Z�Ĩ8�$ A�M�9�o���ګ�VX
q'�@��ASO��7qc���&�<��$��g���2
�i�a"A)p����e�_9�0O�Z�{��ZM豂+	�&���������{�D��0�z�Y�ND�X�K+9�|t`�����C�/��o��rq`�N3�s��!!]��¨,B�,�/t�=3C�r�:��ۢ$h<	�Ƀ	����$nɆ���Ֆ��g�4FJ�Tޖ��t*Ϋ�����ˉYk�K-�� ��۔Э�MZ�5�5*�A[�z���yb�}�K�� �9��ëp�狴�E�p)�<�?��Z��E=�������`BlY㐊E�ح��aK4����-_8v4FB8��j.@���M�K���oJ��rzv Ԅz�`��IgՋ�r7��)Z�$P�����^���}��ܭ�w������D\�9]<�=�yzY�H%6*��XI0i�tqHB��I�jcm˝���.�w�������Ў:j,���k���q��{E�(AZ8�����A?�T�������ɝ��Ob�o�s8�x���Q�Nթ���?cx�>x\���xaT��=2"�v�Y�'��SD˫T�䰢�ReI9�K6�GVS0;�(_
�a�����dEO�?_�˖�'5\�veF�v�20J�>=�Q1;����iMd�v,��
��^�3���{@߸U}�{A�X�ߒ�U�Y�H��m�o��/�p��M��� �z%���޸f�ps}�Y��'��J9@�Kɋ�Ui��zW�|���&#ݜ����Wt��1 ��	��
#R(���i�(��!J�W׭t�Za]W���9��	�Χ��j�(Mh��f�<�g}0��|�1o��5�Gm����+�8�� &��.�<�p��!@���5ԌHW{���!|��!�0�L�6�yBL�c���!�/�T��^d0(�Ŭ�i�W��.��΃9�������"��'���C2o���J�1�-�[jC[�Ӄ�ea������dYN.�Gh�������)�'��;��k�b����W���C�ȥڙ2KEV'O��������Y��<���XB�TW^��6W�\�4�-��!���31R���琢
%S�1�)?��h^�N��(����Tx�U��.��KY�C��8��J�U���]��9#�Ī0�Q���K5��֦��%[�#"�1i���τS�L��>�BsS~'�0�Q܌�����@��F���D����9XKbg����Yė�1��hN��r����M?+�i܅ī�� ��cΓ OF˘>q�j;c�lx�Y����9�~8rJ�Rb,�0b��7'��Cwz�4K&8��}߁lf}P�o�����~��"����
t��/?�%K�I�C�Vל�&7�&�(���7{���a��e���L.u	p����KAW��\.*�-�[�r��d>����q��n�m]�am��L��"f�h��g�����A=��9(V�TR�Te�E�C�n�ԃӏ^r??v�N���wӇr���o��/�����.pu���Ts��:���th��#���!k��q^Dd�����v'cq��;a�u��]��O��.��n���`|�<���ӥ[{�.�q��zwi��%������,I �Pԯm�F�H�3@yn�#�����jG�P�r�'�]��\N�(̃ �?���lm�J^)_�J�6�<����i*��j��K�Ksy�r�(s'��u;&��pz���ki��R�RyKc�$�$�Dت�%�^����;���ȱ���-9�rP]d⍏�>k�Kz��߽�����,S�
�6�X���$�������4^��t�"VM1���G6L��m�{�ꈿ[vz�"֢GS�4
�۞��w��Ud�B�'%��iL"���:.ثQ
	��#<t��߅Y[�(2���xu�e��Dz� ��Ӎ0	O▌NC�;�S[8J�Z]�M�[Ec�('i����Ĝua���k�#����G<>2h[ZG��2�l�|�Of�;�!���c��R�"�B���]��i ��6M%	8�P%0�k�TD��_����Aw
�8���l�i�x������p׸��+�ޙT��.��>[�����&첚yr�\���nC�*��"(��p�H�`N��\��u�i�]Z`z\����!�6��;�+t�t�f�������Tn�~�$A�1H<M5��N���q��?��`@y�N�C���s�j ���.F�O8ٰ�a��ҹ�Ӡ]�ql�3�ο����9T�p���=������S�&/cI����ᚬ����9v���>M����5����=�Jb|(�wYMY�y�tn�r�(9�#H1�A��	���o�0UW���L����|D��<FVxd��r�a�yQ6�X1*�Q3���s��uQ ����0v�� ��$��.���d�Yb��xe�0�W��c�*{���(gW�F�/�ɰ�e1"b!签���Y༤+0T���a��j�zx�q�sUiq���jy� UI� x�M[.6"��5��]��t��p9��h����"O[��N#F��8����hf��]���Q���(T�e�`�Ĭ��Wcv����'X.�*�S��*�����1S�%l���%omjߌk��Q�4�����^�Mл>�震�U�k�Q��1�J��\�����jp)I]>� �7�nzz�Eͷ]E�)�H����Ļȅ�dB��E�IFT3�XD��vc,���T~��0q.^�&N_F?r�ې��Ww��ox&��W)}L�<�k�(�T����_Ff�;�f�/R�[ݥm�}~}bA�D5���ԛ��Kr5���
ȱ����̟�]�(nQɮp�B�y\��m�ƈ�q:�(�S��f`�I �g�Y�s�^n6���g�������WH��2v�n�I�^l�,��yĴ���고��f��a�BU�� ���J8��esq�qt���ǂ��������}�	v�Q�C+�7*�� ���}H��0��.*G��'%r`��B8E~����׽������]�g2���?d��l���|�� ��i��\~�p���I� O�8k9J�<p�t�)��8w��U ���%^{XԼq�UPͷ^YY4�E����M[Ϊ(3�z�|A5������IL��~�K�{��ȧH�� �����*�ٚͶ�M�W�{�5`(f���ڣ���ׁ�*ݝH���B�Ns����?�6qT&�����a#�	kS�������U�%�\�H��C��퀜���̠��k��>�)��@=e��V�����W�m�Fǈ�T��[ʇv9�Ԥ �W=�b#b��[>����Pg�7�+A~#�Ź�Qi�ZyH����i���e������%��e�$|T3-�`�o	��3b!�I:�s���ր�bF���4ʜ�|�ƱBa�}O?n�Y0���z���tT���bZ}�����0,���*���NPu����	����$�M��Vx(����m�vׅ�dI�?<')��n�݆{�#5>yu��Aqw�ecc��%(w���'��A86Z㔣@�롴ŭ챹t/({�G��X25�����i���T����������tϱ�̑��u��)��8��� �"
�N��މ��ݧSqq�%t�i�D�0�ڂ��`�_y�7ԓv��-�s>eM.��8(�zo�6��Y�IL�?������k�z�{�]�q��PY�z��e׉��^�q�����Ⱥ���yo�8`�_B>]ѩ
�=P���k�'�unp^���5\KS��=��t}��ړ¼k���݅ͮ	>Έ��K��H�I�w�,�q�����e�)�l�Ű�w`b����bϭ�+��g �T9��ݮ*A�M/
ɏ�%��7���KH/w;u��Q^T. T�z�yS�F��͈�w��?Z|CH�+��2S΁(��y�v�����7�[ٹ� �M�[�~�O��ޔ��M���\u���Č���[Q>���a�R=�5ӎ>�x�p���_�tx�ia�|��������!b5�_8ޕ����"���a���N�G߮r�Q�]�7U.��l%\���$?4�N_v�-6<Q8i|G�4h�TQc�8����Ս[�ֆ6�_z��3d>!;�>z<�Mz����2�%���v�=�Χ ���(��;�LD�L��h�R�p���� ���*��"��/or���b����:��UR�����Z��O���w����R����wew�:oUy8���sC��b�,O�|�+֘���Z7�a�<я��>N�����|T��y���ap&E�1�BI�~��,���a6ÍU/Z�s�Q���n�u��
�|���:7P�]��1{M��1T�=/Q+���_��CZ'�Y^�>�?0"���w�4�O�xJ藮0λ����k�K�1������-��T�Ae�F�GFĳ�ˍ��&:5����v��[gg���Ptڷ�;�������}�)�4�hD��:�8d���'vA���}��Ȓ#�,�7�!?��GG��w�@�`Z�ŵۺ�!:���k2���m�����v�_�3���,���V_{��t�{VҲ%h�p��Ǵ�O"�c�.���cF� �=��mIE�޸k�O�ɁR�
�@|�)����G�0�x�K�&�]c���S��D7�2��N�����Tu�����5�sַ����&}n�/�P��"I��>��J��L��>s�+�X~RK�]Vë���>�y}G��G����q%Ճk���p����9{���Y����K�ǃLJ���x���㞮���C��S�[�$B�;�'�sc�ϟ������̧Ge/����t�E��9�{���1��g��EOU�ܺu��W��؎�\Z}
U�On�T:Aذ�����ɨ��r�c���������;4x��?���h_��Y�2����. ˜?f�^l�VsmI��ۡ� ��;�?e��j��gm�����,�"Nk�ZC�㖹�B������6��0W�?S�g��L�>�� &}�\-7�����(����7c��;m7Z�!����M�#E�T���$@-dg�7dn|�K7��#N���q�������g̕��v�'��d��Qg����������Ñ�e�Ѻ�.��r�H=t䟢E���м#���q��D���ŕ�.Zs�׏��.�gUm�?��;)x���骧ǿ�PС�'��������o<��:�y|}
��v��1�ŘU�5���]���N� ��$� �"���H��r�a5��ǫ�^/}��:r�,}.�.tX �bP��Q6��"�Z�Ǟ��O��V��kՁ#|@���q� ��G�1~����3���S�����~���J�8g�w��{Τ����H���t���o���1R�}bf��7��*�H�-��k(=�#�>�\����R���H�������]�,u-�P�;��Nj9����v}{�R�=���:-�_C��^39����D��^����?�rT93����
���S<���zn����#y��[m�4(�A�3�DsH�@P�#C��O4gG��N`\!f�Wӟ��b8Q"#�"�e�ؗ6�Y\�������1k�i�_��oH����6Iќ�\y��SK��':w����>�*H� VL�7�,cq��?�ų�p]Ra��D��xi��Y������_u�b��~���#�t�r���Ma	�\����n��^���*hM.�=��0,�W440�%J�x��;1��-Wy���<m�����j�|C��E���l���\��:������wzݍ*=,"ҵSٺ�v�Һ��W,&xb���A9��k��c�Q֣��S�S���	A �<u�XW}�;�����X���Ek��ȴ�K��S�TV���'e_"��/�R˵o[�C�+�pAs�gba�x��]�/%��!c��^\ǌ'Q矸�i̜���!���=RSU\���2�R�\�9�T>���ߞ�Z���a^MC����j���>a�Ã�ŭA�'3��3L�򀴓�߄�ٸW1da�O�_���F�����3P��_�~u���R8ak��ZWnm&;�.�w����X�����Y_)LP��	��k�{e�nH���&�B����xJ���T�~P�#��q��S�S�<m�5i�qv$��ק���Պ�PH�J���sc���U�$��%�5��y�:�^��K�|*��7*�����ֲ�g�JK]��v+x*5�вl-	Gt��Uש��*��K�e�L������r�]w
1R1*��?�yb$vp8 *	u��5�	�L��(	bF����P�."��k&?N�4<q"�2�w�D��ͮR�$�w���ʳ#л� Cv��~)���d�جy vj���ņ�`V��K_Oj=q���}��M;��粔��eP��l�bTds�Z4;f���9���6�h�;S�^�5��X?'�N�IE\H�HϪv�s����4޺�cM�{V�:�q=�
�O��r�>���g�B�B=Y5�#)������n�4	&� e���UW�+sLn{$��v~h��Z�/��(�ᳶb�,����3H	�<�)�.�{��e�����M�iZ����$�j"ً����ol<�Z�%\�����%�_�����GC�NL��2T��(&�|(aG�[�V����;�����E�D��]��@� H��u�ʱ+V�	�|��t-+�����[[ۜ�:����y�E�F3?ٍK-2]E�Ҽ�#�̾��s6��6��DIY/Χ��o�]Ag%��	�(��5�T�Z�+V;��˚{�X׀��b�c��T/�RH0�t��˅9�+��dm+�@�46Z��ц�Hz��h�V��2�9;=7=����T�F}�JLd�ɨ�P{����M�+2�j�dw&2q�ڼ�ZS2��@��M9�LX�
��9�����!u��Ov���j�%�sM*����@=��Ft�fB��X�t��6�����2R\�L�a�_yl���__"�K��nm_c$D;���(�B��,�i�rM2r-����ދys�gQB�H�r��b�JG��,ia�:�Q��mw��]��㥐������G�� ���� F����k%	�ф�}���0���P�W8|c_� (��eI"�0npL@�吵(Y�^��m�7ܝqY�YK��hF�΀���S�5������%ӄ��p�S}%��������0aQ�3*������%c������oCI�и�����tw�b׸�Ԉ��d�y���Z�aD��&O�&�#��Vzn�T�F�FT�-h���a��9�ξD�͟��Sw	����үq�icu�_ iŞ!WC��Z뷩�3�r@^8��R���q�[��?n���|��P�/L|`/�����bj�^%ڜC]q�
nl����jM�VoG������-l҂t�H�ͶO�_'<�cj�F6_��T��珮s5��.��A�!]��J��m������̨+iKJ��MO\~y_Y��"!���kTZV�zZjj��5}!%曇�w�9k��J}�ۑ�t�0�j�WU�\��I�R�Ҡ�K���:�2݆��$���^ʭ����y��8.���u:[@�f��p�׬��]�F��t���s}��n;���p�<���H����6^k
�>
<���sg�/��ϵ��Hy��4q�R�&�♬O\�a�UsZ��X�O���T�D�A�#0Gq�S�F��Ћ��=�L.��8�L�VY���Lζ횞�@�{5_�FFa#7u���chSO�V��>����w w"�,NF��,j��??`�
Z��+;51�I���/o���:�v�����{P��\�n��9�62��~2��{	"�;�oPh��)�[�C�����H�Z�!m`�G<�uL:�����Fc���ɡ����ɩ�_�)e� Qm��D��ʡ"p���X:|��5��
�!QߙQ��(!>���&�Q�gQs����4���	���H�㢺���۾��A��s�>&�_`<O��(B;�i��ݡ�<�51�I��W��=�ڎk]Ea'0n&$km�#���Օ��Aas#��˽\�2deH���X�I����:9�^�֠���UV?c)�;�"�`�5.�+�][����-x)�]۹������y.���L,D~+L�O����C��.۝E��@R�o�Y��7>A!�5��*R�((���Cٗ�L�� �k*��I�>�-C`n�酋�0��v@�	��R�����1+}s�G3O�Lt�7ȹ�4M뜷i�J�����{G5��}�x8����"�
(M����T�JB�5B�MS�J��"5��IUj�5�P�IHB��.�>[e�q�_w|�{�x�p8�bΧͧ���5�2�+��Lhka�G�t}Z.E�B��r�iw:�S0,�Hs3�� �������z+���y~�2ݪ�ńЛ��?V1o	�k�����֙���h8���8������>`B�})��H.�L"%��sS�l���U��}̪����k+�V���L��<����6�k!��|���߰��˅�=$ο\�k�Qf����$�J��4[���~ԟ8��Q�~2�/=�U�B�I��/�E̩�����!�LA�:)�~�-��% ��$�q�i?M-���iU9���S�ʑbb�1��'�#�2l uFś��K�{��K]N��H������4!��i���rq�-ȯ͆d�����^��0t=����p~K)�W B1\
q�t����'�>#�z�(H@ҏ/-�a�X��㆜c(����]�u�'���$�d�l����A@O�D�!�ȳ�)P�ӳDw��O�
4k I^��mј���Ǘ�(�1�ڏ���H(�d����'�������c;�r/"U��Z��׮ȃb����9��u,3�Ғ�N�pb��`"B�%B.!(q��h�i�%!����O=�q��P�P�#�^�}/���@}`��F�bM��8�*�s���Hi��e���N-qT�v�ke.5�y|H�{���見�4�G�};v�`�c�Y�Xh�BJ6B�p�;
�>a�	&?׳kP�=(UI�+�뫐���<�V><��\G�q딬�Ʋk5�nT�E��^)�e�|�9L88��q{ލ���}~B�̫M��Ő����i�}$T�\�0ݐ��/�0�l�M����Kopu}�\��f\�%��e�J�/�d��!����Я�,7:�!$"��nD�'��Y���>�*���Aγ���{�T�A*FL�@��x@C��-������Đ��N_/3Bd!�F��8 �0�ϩ׷�is�&�Gw��,>�����k�1��K-��{��r^��0��l��Y���2��g��|�t��������w$s�~�%�׫'�>w%���?椈�技�O��\����v�9Un%ÅC�7�=m����.]��l�1��W���6rM`h�( z��XQn�j�JM킑5i7<�	�$xw�&���.F��Џ$V��5�y
0�Do�j��}P��ĺ�J���IXcJ��n:N+��B�OTx-4�r�3VD�>1��J��n�Cm�Ł�X��*݄ �+i�,���X�b��1&S�wj�u� }�H̙=���o�����,�op�kk/=�x,U{�r���u<�	�= ��Z�^���4B�zRX��tE�*{ֹ�־�jKdAp2?đ���Voϰx�X�{e��y�����X���Hg.\���2��rc��GL�kx����)��Z�^b�_�M}k���,�RW�@����w$I�w���:
��J<F����%��HV��6���Q�:���A�쯭Sq)Pbi��@3_:`�Ur����K�)�ɘ�^ݖ���DK�VH9JO��h�q"@�5�QFU�N��>����Ϳ��&w<r�vV�T�D��%�D�قFҧ�\�h��o���������,AZ"��qM����g���M��mv)]Ũ|��ϋ�>����a.�����ģ*X�rl0��1�=K�D:�t�od&8�CFhq���V��GS2�)�!$ޟU��w���-�m��V%Pov�=!��g۾�=�Sb�p�u[��e�[� �I���E��Ab:�F�Jw�������ĬI���ӆ+x �ĵ��UNv��3����k3�l�I�)ʜ�;F��P�lEhåX~��+�h'� ە?�w|�X�j���
m��2o�K��}�|k)��=�/'�Ww8���/�`9��i���W��[q���5#�? 9��: OL�Ǥ~#�:"Z��J��L����鍫�J]����M\D�m�[�þ������a�
���ɛpfs"V��{�[�!B�G�q�i�!� �{�)l7��vc��%�)����I�__�[[}�m|)r_ze׹W��F=�p�����Bׅ�!��<����a�|Jc��`�͗%�ʼ�߫wWY�mm�)
� "�-����H!�v�	lS~�Ǘ��[�!%����5��ƥ���T%C��+�؟�"u,v���Щ ���C�!�G���ī���Xv=�,R���aP�D�����A�	
/G�=�)|ֿ���.�v��e���~h��  ��P�+����bto�f����߂�j�ku\S�gT{K�v�nv�C�v^`5U�1�V�D��zX�!��EW?�FEh
-�E���\&Ѿ_^�&Ͼ��	}�?ɾ������<���D�<JR�z�+.;��k��m��E�/V�5����p
���˯/���@� ���%�ǜ�Z	�e��a��+���.����? gM����/ u�=��s�� ����4����������Ə�_�J��M?�F⺭$DS��'��ѡC�ſ��M���㛳�e�U	g2
z�h�K�g�� ����n�\���Wg����;cdd��XM�u�a�z�F�ֱ�o�9�Y9�ԡ��2J|4&ꎎPI�?��Cq@aD�7 ��������Եoov5����y�YͲ�&�)zW�LW��p~���A��g}�?;�7�	e��ubK��t3�ht!�r�oh �d���Θkq+��?�zY;�UZ��&��%,l�g�5's8�b�Qߘ���3:���"mʭ��oQ ��ugߑ��X�b
�߹i�����<�ϥ(�E)�ͻ�Y���F0��1~U{êaB	e���� @󜫋�cJ��Jl`vW]����X)W�M�moۚ���Ur[��Іq�������7!������.��k����'�� ���r�sHX_�?; `�K���I>��ߞ�I~�w|4f3Af�С���3t7�H?�������Z�-tJU^���:%
u�I;`�eZ�ǘ�13k�5�!�-Z�������B���GI�^{;�Z���e`5�
r����~�e��Y�2}�|��r`樯҄�孬\�Ǒs�su<�RTT���4h���~î<1
a�X'u��Zt0��گy1��%�s\5���Dw� s%F%�}�����,_���򾾸��r������:Q�U��\v�	?�zm(�s��m�Lze�� ��<�Y�l$�09N<�rZvA�򓚧&�mr	�]op����ؖ����),������3G{��u^�Ǿ#ߒ�j�Ȉ�(�UءWO�ϟ�ZިU�Z���,���s����d�s1��G����3��~j^dR������H�٩�:���3$ރ��9^��3 ��^�;v�vN�d��*��|ǛB$ħ��V@,9g�vf�ZP���+jNx������;9V�>�k����B�7�w�(bC� �L/	�c��f��D!��98Ny��!Hʢ_�C�s�t�@5rl\�26JU�$��`c��C���G�d���f&5�`1&��9��� �(hw����@���P*lnh{�J��vz9̫%У����K���������T������Vf*�hY���]�7OZ���Qt��IØ��G�;�vƈ�m`�ȷ�7|=:���/�My������(w�jώ�6�: ��`�6=q����g�����v��[�9_<Ro2Q�*v4s�
�e-��[Ԏ��Gk��K��w�(A�G�||�d�<���6ޏ��T0��iZS�7l�����t#i�s㾵�I�9Tb�qG��[�|M�N�p�~*׹�����kY�p�p5FК��#��xj&*�z��~Y�Lv�ȍ�铐�ҳ�!P�B�k�fZ�k�`� �a*T�E� Ewٔ�f���s.�P"�t�
�����������%��qG�j�;�'&q��a��^	2���TR��I @���m7�M�W۞
�`�wA��ϱe�X�g#|���ے+�%^+���KqF�@�ʳԒ������w?�ׄ��{پ�z�>w�ԏ���'j��C����;�B@Q�J׃͎<Y��P��r�}��{�����ψ��7�B�����qɧ~a�@�R��m� �羠��.9��6���v[���h�C�P��_��0��"�M�{�e*#/�W�e��
k1��Rz��y�E�G�S���p�(�Y��x,CIK���!���.�]߫�o�|�3 &7�f#�SD�Wm��ܶ��E!F����� �K�il���#9��|�n�f,�N���s�����y~^���->k⬍����u�o���A���ͯX�*A^Xo�L%�,������%y����:-�F0�F�3oH��X ގu��q���e�Q����O��������HD��_) ��>�X�}�aO����3{�ݘ�E=�4��0�T;�`��y��o�YՃP����è�7vf��^9����5m��i$�?����`�Vj���z�@%a��=�c����Fq�:[?�2�m�x[s]�}����[����
7�����D!=�oب�^+%���=B-Wעӫ�쇫$-"�\	�Jb��1�o��0�1߶W�z	b�q�f��G[�1f��i(�s'I�/}��� Yp���j� gnÓZ�<wG%���X��+/��I��'��bv�H�����y�ԁu�:�$��硙��/}��Dݝ�ӍeN;�WFi��D�!}�@.UA}/�Q�_��{_��������� ��Q����8��m����b��Dַ8��M�Z4ql�o��.��-�����Ę���sM�����՗,3��{;�n�W.U��ۑ�%����"M��H`F�4�&׿m����r(JP�PK�� 8�X:�ߠ���m�v��Ό �� w�"��Z9'3(p�sW1�`x_A��z�z�z]�@��v�k��f7�����Ef�ʚ�^S:��8*�?%~0h&��eos�d4�=�A���5GOmKXT~���Z�VJ�ɍ�u]��cq��v?ہ��`�(��@g��ɯ]�H��8P���C�}{*|�ѹ�(u�?!l���R�K��3���ȁ��L*w?�6�<\�����ԓ�'P�1$��l��5&�a=H�XmPW�o{v6�66���g\0dаj�ݬ�PCŃK��j���' ]3�c5�}�Pe�����Wt�1<���F���p�=y�x�´�ka�����l߷T_r�Ha
��r<h�f��x�3㿙/�M܇�@9�vV�f�n�%��:����>gl��xAc�����Q=ح21s�-F䚀jy�U7!͏ˍ���5����P2oP�X�w5q_֢ɞ!!�(3�	�\��|�,#F�W���t���0٭)�mI�k�t�o�",�aDLU|z�����1��¹F���Ċ�w岲�E	��9��{�IdP�( �GS3�V.`�X�����>leD֤\IІg���e�4X�������\LZ��e<F�7�c��7
f݅�,4K�btg�Z�|p�e�a�ֻ�tA�~�3���N�������7��q8:i��Aa*vS_���t\OO
�,.z��tg���
��2��f����;%����n ���pۿ��3���	�mD��׃Z&�*��%�ԛ�a�)̐��EKgB�J~yAy�%��
���w~B�$]��N z�e���M�x�7L0���P.$�sI�H�Ȍ���B�D��[k��6�x��U�/�|i�X�E��0����r���@t[��|+� ?�#����&��Z�yZ�ȨE�fx�.f���n��`7E�ѱo�� `&T(C�fg-Bls=[��nvx��w]�|n���d`�@��xbl����~E��u�r�M(,V)Nk�����a���a,�5���,7o�!��E;�����c���&�Ҫ2kX<�G��X�/qR�͇{-K�*�E�Y�2^��f���@ݔ"O��cW>�r$�h7�{|n��R|+"MŠ��w��'�Dyz��L�\����^��U���"�p�"z�a��9��ӳda�s��m���#Q������78�؍�@��{a{����\A�p#�=�<u�SKQ]�:����v�����F����0�]�]��F{�����t������A�z�(w�i9jj��?x�p�yY�]�~�b�nL��ꋷ�����|�s�5��Uܱ�5�w,�8��`�x "� 6����O��<�]��f�`�ePa�֛gP��k%u�7�����'�@�5��.��rE�De0�������`��X1�#���KkK�d���U��N�*�՝f_R�蒁nvc�1S�Q�+/�6IǷ�~���ߠ>��#��O�������v�E��{ZH�,7�1�s����|�mt�:���!�(?�%��U��lpe��V+��S�I�ΐF�A�=ʱ��o�6j?�O��~,���mbu�s�W���+$հ�JQ�ff��'���|;{5�ّj,w��s�f	�����G��ט�qN�Ǉj�v��.8��<B�|�y �����t�K����jnv���U�� v2��z�z����Kx���i.|�Whm�.�����rFv2L���4x��a��N2�!�8�Q���Χj��#��u>U f�Y�N��+,%O`�sJ��Ŀm�,��6v��")Ö�g�'���`��}�KM�^" |
����b_ly�困1R;,��V��Wk���<�a�D��᠊T���V:&(ѣ�������d���1VD=^c1��ȣ�fKH��E� ��X�JFVڔU~ed��En��8r.DH������B�� L��$��خԿeV_��h?�E�ت�[Z�2go��n$�L��b�$+3���4�[�2[�;�� 2��"�K�Ap��%Խ�b�l��ÆGv�C�U�]�A���U��@�Z]��ӔD�����pWt�5���j*J�6GL��aZ|���R�ĸrI�w�.	|d{���G�JKyI�Fm.�\�b^�J���ռ� m����W����4��	����o�וP&D]9�h��h�~�޽����0�L�
Y���n�2�uwB؝���u9B����2fI���b�x���8���%��B�ƌ���*d7���z�H@��C�� � �M}������i�x*}/�*X�W�0o�*>�:�C�b����Q�{��(��	�XF�d�_��ٳz�jя�2:�^�b�N�x�n�NeYAU�~2+����z�c�`3���d�{�L��դM�a΀-����f|�2���yij���M���I�sI�
>^ݾ�a~��Tu���`�ࠥT*'��ϠL/����Ȉ:��y^�P���ያ�������ݟl�?̒�E�>�צEVy<�^�VGe�)w��/v?���0����	�M@p{��PW#�Ƅ4�9�TO�t�;�Dq9��{��ñc�����v�ug��*7Zڀ��*���<���IV�nq�be��;�ߝݬ$��y[�d��lT%���Ae��W}�ׄ��f���]�<G-:}�e+�����A��,��f�$N��QK0ǭ��C�3#@}&8���~��´�5Ş\� ��ڃJ@�(?Ѓ��_��p��"LBc� �&yh���qfpCQ	�C ���F��P�{�xk�,��\&�
B�2�N�cJ䫎��M�-��x!�)�P�i����E�C���[>H��^��j8���"������Cc��&���yr�?Pm��[�gH]���a��!3pąBN  �E�H�?H����������S̠���s:ˆ�UX���J�~�6��|nJ^�=�z�PEQ5�a���&vw���0�|��z%�
��p���&t���r��am��ܚ�J�iGγ�
1`�j�!�T��j0����#�\��o�Z�!�vD�>?���Jry��kY
�4@XwD{��6��g��-���>�i7ZO�+?HM�������������Y7J�F�Tuv��0�҅x T��-l,|�Nb���؄�����|ܵ��1P���+*������_�N���[KW�X��/"7la'�%hh�}-`��.�С�\�x[u��.j��`��*�~�ldɖ�wp05ȭ�9��[��"�N�Nu:�e���ݕ��=�6(U;������5��.��B��N� Ƈ+��X|���ee�8�
F�����.��<kNRG^���"�|�m���6�I�>���%�l����T���k���g�d��OI�ɇKK���I��o{s@�G�]$����-������u�rӲ#���j"����_f�C�9�
$�_**���o@ɺ��+	�ꂔ�v��I�g��u��oP�2��(�;F�%lxmϖj�a�v�78��1�,�E�����d�����.D�4*H�m�Ԁ��K��s�c#��*a��)�<�Iɢ���B�,�.���͐!F����5gB�Kx��-��s�ZZ�Z4�K����R⹊��\�L�X^�7�PFA�V�''USY��VRp�՛����R�������{S;���w�[v��	8o4�8�	�8�L��g���2�{��:袌o�M�E�a�TH��d������%�5o���r�,�7��7=\O��PFC-�Jb�t��\�NC�e�`�/��>��M�HiL$]vf���p	�={�T�2�b�8�)9E�+2w��.���"��ē��>6q�C�=���59̐��7/�����Z�88���v���C.�N�:y�����VwN��9y6����2�O���_���2�q��#�R]?����ڙK��u�������-4�k,c6q�cN�Q�;���k�Bh�`�:�	Q��8n���JO#/���ɧ��G�Pr����=b�����`?������P}i!��m/m+X���vN��|����]qU����.�L�'T/˜R-�N�����p"�u��9�S:�A)�#I��9J����]�7 rE�����!ɧ�
U}F�R���"瞛S�3���!ԇ��A8���.Fh���Ј��;�9�T_��XN8��\����,��ꤖ��$�eI�J���`���؟e��[<��O��)��eh�m��e*#�\���J-�ow\6���@O0{k7�_�Z��{�
j��o)"�'Ѵ�?�#��r�( ����:��ȤW�0o{��DNQ(!|y�{~)�9PhB�C�,}Xp+��0cQ����ܱ`���X�цH�jNHSa;1�6V%��6k�\�0ޚ��0#/'L��_
O~�k�y�+��M�� r�˂��-�۔�ڼ[+��@>X��be�E1x�{����s�@�O�?��m����U�:<� ���h����24��[���I�q�;�c�ߐ��He�>�c��J�E���ꇵ}9�ǹ���e�HS�e�)'�W�`��a!����Ӣ6�`�ߵ6��!���2���'m��!����u mf%M��&|6����˛ o�r#�qrBE�!�u�� �j-����/|t��q��׎����a���$y|��BW�n����v�����;J�\�@�v�i����{������]S�R��X��K����s�Boȿ�*��p�,�hP����c7LDP$�����\���:V�-MPK�F��x��Ѓ��;��^�G���o��Ei�� '����CKXr�Z��0��p�����`"pb<�HuK��`�a:�5�fT�p�d1��wU'���U�8|
l:��;!�!��'����o�����2�_���1}���wH9�+�����fnBwA�v��VE������+Ayjv�D"�<i�4�З)��X�.�`���y&ݖ��Nz~����=܀�#r����q-[}���[=.�	���	ư����8	�~��tvH��30��m�jy�R����ك����Z����.�4����"g�Y���d���&��-��Vğ��li��$��S,� )�,^�.�eG���
q���3`�*�x�,7�c�"' ��@�k� NZ�.�<~`*��W�Z)�Li<H���܇6��MB��%�J�s������������,D�>��-��I��Ʒ������K	5o�k�+�:�I����sKo�Q�3m���z�F �����>Je��||k�����Q�E����\�E�h�Le�z�a�M��2,Ë�ɳ��: ��t��п1 P����0�œ����+���9��{�SAF^"@�t 
=���AV�� PF��ȏ���K�X���1�3Z�q���obqg�.�5,�".YU���^H���
0���O���e̹L��V�mu6�-��&�Y����f���NM�_.�?-Ks��W�\��,�����9e��$d5t�Il/lxb��3��Z�>/�<��.�����տl�ff�n��S~��}v��Gå�9fN�;�2F�'ࢌ��,_�[}J�<�)�Ex��PT��1�9��]G���H�|�9𧞳zx�?�B+Gw�ɡ#;��:�Ò�V���l�s�k��~�oN|�ҁ$��uGȋ���cdŅ���$v���B:���J�|���*���j�[,�^�fߺ��vL��=�i���1?���ඵ��>s	L��E���������=�ҍ�G��a���!��2,�7\�#��^z4�7�`�+D��6�"���� ���#��23�}��(���0L�c�/I��ga22���w�?�-�~��G��߃'����c��1�Ӽ}�f��뎙��}�o(3�[������:A�!d �#�,s�+���jy�q�������.�Y�R�PMPJM�3�j~��6��u)v��~��?��IBw���۞�9��]���7��)!��z�]I9
�WF0�g~���� �ph麱� ��l Ud�ų���D����S������e����a��-7�m8:��Ǽ�R���&Fs���Z��i3��ܠ��&�ԓ�\�g�zճƲp�v��n��E?>�Q!?1��3}�ApSg�� 7Y7j�8���Ym"��9�1�f���1(�Y�{�c���IG�]�GyI9��FN1�b+">�m�J�i�����G6\y<�w�x����|7�16f�]bҧ �?����� �sb�o9<�G�Y�m��(�Y���Gx�<��0?���~w�J$�u���۾?���� �+O�|�-��
�^ѣ3��f�M �[����3ԦN�(���������8|����_uj�Y���b�B��8�-\Q�wM��ZNԉYd�f��`���Oc��C�R3�o��9��P�34� L�NL{��1��N���˧SF�r0�jS����Z�f�Q	1J����ӤY��)f�z_�jd�q833�[�q�X�#'M�Kl�ع�/�y3Nk#:;��\&�M
���6�6?z��G�o�I;�Ƅ�ό �Ԭ����u8E����}̉��-�I������V����^h'�i�AĒ�n2�C���m�;�y��~�jn�O̒~���s��g<�s�ɢ9T)>��J5�g~��r.�r£^��\0�t�Z��E��r_w��-�2�(NPW��Ihϲ���-�,��Z����-g�
]����@]����>݉f`��D��oc�H�٭�s$2}�).�o�\_����C�����E����1�z��P�;���WO��M;0�̶
 p�e>`�*T���,R5̔8��s�XT��3����A���A��?��� �~�s;b��p�6�!��4+����V��9pG �Q3��h�:ԧ*����eD���412���?Vu/]��6r:�BW3�/�~o�` s� ĸ@�f��(�L����8�lՑ��U�1m��6[[?	ׯg81α=C[�=��瀜tڃ����rN�����o	$�]���|gX�QT��ۙ�*+g���9π��ׁ�=���g���/v2��}U	�y�|@������M��:v���?���y�����S� ֤S�����4��"���5�6�sN%��Gs�y�6��O����n���V�|9N�����7��TT�t�����7�F���%���V��������xEsV����z$ne�L0q������@�i�U��9W������^ssv.�?���H���V�9�B��h�C:n�����=5�,^7�n'���>H�>�V�U�_sd�W@���E�\Wqk�9��jh��7{������aq�g���#�e<-�x�#������;��5@�@���l_r�O������s6#�[	LΗu{oi5���W>��S�/#�P�G:C���)=P印{*c�`O�b��������+9DgC��;�HX��q�e;\�����=��a�9���\t��ZC�!l)c�_�K��^���<����V��Ay����}�\���05��F�*{�x��3���]�](���27
�_�lgvL
���,.�y�
��>R.x��5k] B���(i/y��B���7�T�J�T���E�X�D�X2z�O���
��I�5�I�7{���Żo��z1��A�sa�<A�-sH���d��!2%�}�L,X`�uż��{��q�����a����AAT��ƅ6���b���<Y�Ve�WJ)5��>G=�6��0�gl��::�J��-5�;G���f��X�e�)���|��`��r���<���O���%�W��H���,���R���	�|��MS_h��/$">�s䲰�.eFݙ�5jOd/ó]��|���Ա/>�7��h��5���k�e"�U�� �	��ѩsZ�jiF��|b zڷ`_���.+����+�*�H�]s��?��]]�,8q;��M�,#ڌP�3�8�l��x��x?��A�j��T�]�\���0���2��ގ�3���]���G�^���7���o�%>O�y��W��,O�����l��IQ��\�n�ս���t6��0����^G4R{�*gJv�[	�9�⇢��g`�����ބ�-��D�E=��%����t�����ܼ����f�F�ͮi!�^+ݽ��m3u�2{���t(�A2�7c�y%�|ߌ&r�Bu�x�8:�ù�L�D����֤���v׏q��=��"��a�8[��msW�:����\5Q�{]�_�>er V�}�)�5toSn���@�������axP�P�����Q���*QR���P?#!���3���챭����ѷ?���qQ�}s����,���Y�|A�:5����D?�Hfǀ�Mn���0md��G�������Y����٠�m�4�-O��94�n~q"���;zg!�1�'��:ccA=`��W����4\�@����5��\�=��A����çxUX���ۮiO��������,?�������Ѣ�nfw�`a��rU�}&V�fȵ����[�aGQRE�g_�쎞����4L����O֒�-%��G�Dҧ��T������@cq��z��¢C���v�)���\ԕ����t�F�zp�����C�F�Գ�Y����o?����?�Q<�p�g� $�+vwr܁R[�����QtS��X��Te�����*�ǤӃ���������mB�G�v�UQ�oD�'5���߫5r5U[��H@�+_�0��iTxv�7��<'�s����Z%��X����t}=�S79�R��(XB�e�d�@b{̮x.�\м&CF6���K�)a�QĽ)�o5�4荊j���7-	hV�dݣT����s��*�;��$���h�=�lߨ�;�e!�c�G�u�Kmm`�2�����i�yA<lb�]<i�+�W��m���.}D�{��,k�O�P�����KU�S���Fu���u�{�h��MN3��M��k�1����E�F�$��MH������id�zV6%�<�s������^���8m��OV�{��h�\�)4-NXN��=���}��������u/�\�x�Q9�#h��J�5)�!�'�!�)ˮ�3�A4Qoz�f�sL�6����oՔB�b;�Έ#�=�Û�zLw5�>?&(4�A����t������&�"�#E�"����0�+�����j ��3�$��U���)ݠ���]ž��¬Uȕ��>�}���.��?&??���KAC2DL 2��r�qkt$���7�;	���n5�F��J���V�6��:�-���K�U|L��s`c֘6n;{��Ln�\����vK�4��r=��"���=�Q�@@���^�+@����HT�aa��[����8qkl$�1����-2�u8['�ͧ����Fը8�tH;-�
[��G��v�U}#�7�"g���̣:�>��7ne�߻�ݞ�o6 �D���`v2=��MR�g
�}}r�u�T�4�Q�ܐ����dE�d�;}!�\�@�<��c��5?��Q���.ٻﱜ7����Rq<ҳٴ�ʟ6X���T�Z������I�ln�����w�r��	+��֕M."�~P��i1&�������Ӊ&j�Y{�B�\���C$��{���kq�_���UG��!�L�Qå��e��4�+��Yfژ��?<V��H�L[�cO�D��
D_o�P)��Z�C�dʭŖ�6�tRB��2܁֘E�qv��s��_lVU��ya�ȵ��I�����SI�zڕ,~yB+G�?���7A�3�}�M�(��`��1�)�$G��.K(�x���)���6�n�,4�(�o��b����I�5�m���N� ��"<�F�S�>])i�o�t�[ׂ��P';�ڛ��׫$���b���L�zcr����D��>�;ZœP7M�Y$8����`��Q�����n=�X��6���Ou�����^�?J��;���(�7w�%}��l4˯������D�ؙ��_���5�����^�?ub�H��恷��'}7�Ԓ��P��W�_��)"^V��-�1O�	d��^Myc�ʫ'��-�f���P�M�ta��'g��\���g�J�j���Dt{� M���R����E��v��� 6O���Q���y|�Z���q�i���n]W�f�X�;�k�Ş�S8c0��h�Ƙ8Jnq� �]�f���L��q((y%E��~�������P�n�hda8ŉi@���\��V���Z;s���(q�P����h�|nX2�\�F[AT��D�M�2�W�����Q��N���!������5�@�(j�u�g)�+y�6��A�ϒ�i
³I���u�ZDU&�l��$D������Y�g[�R�A���^@�|��C/G���zH
�}~�FmH�����+/�oܺE����C��w��߸z-,�M}�S#W#=�����w2���` �Yp�H�>�������U~(�4JH�T��CV�>7>��N;�v��JZ&-W���b��di��}U��׿S���*%���Z5��6�y�TKEf�R���\�Q���~�披t���
�kK5e+���8��3��Awe��=J��Ǝ���/uJ��.�����=ݲ��C �r�ny�g���<����5��vO4�wt`T6J�ǂg�܆�TZ]�N�ܯ/Cղ�ق��m��)�,�����R��r�l�u7�L�M��z�_���Ww�n�y>qS4���-�J��y�
q�g��L#���f����X��,�f��I۸k������9m�ʉ"�W�J����q�x��&4:}Y���>�ܩ���B������3>���z��������`� D#���r�l�B���f'(���C̈��֪����u�ud�ɭ�sp>4��F�S�wH�0��5:ELq�;��]������!�Ç�[ ������
�f�!/*�O:��O��w�>kԒ&Fa�/���(��o��#����������:z��<+3S�����b5_��vds"�>��]ͷ`�Ʃ���sa��d��4˥��@��y��e}z�Ґw�N���z�F��y�rx�Q%��O&�����Z�ph�B��3&��5v�Βq����__�(:
+1N���I>Z�ҀNv�����8��A��b ��Fm��N�v ����3�[�+}��,�z�Q�?++�\���^cs�r�<a�%~l�;�E��� wr5OM�� �(�a�D��B�{��@_6���`p[5�9 �tK��-9�ԚJ	(I~� [b���4fN�m>����^����9�9���]?�Di�*���a2I[G�����m,=���	�t��9����7y�k�,^ӓ�K�.���i�&q�^yxj&]E�u��+>r����7��'uR ���+�c�}�/��
���eW�?"l�c<7'�7ߊ.(ڈ���+B[��vOcP#��,��k��R�,e�(��УU�L�ۖr&��(Uk	C+~���E�{�ad-��Ks�������������e^�ioi� ��Ro���G�ѕ�,̕Z��P��n]�=�oeq�Xm��mJ��j�ՄN��v�/>νa/ΰȫ�|�ᧀ0��M�V6�6{���t�("l��q��(������M{o�l���2���>+#K!���8���d�v-�kp����실�/饸N�"5�ՖZo��N�i�J�\���!��פߐ��=�QG�K >�VHR:�@T����(�#sy��䴥��������� --b�����tV��4���_�ϱ�nC��9�9���͍�Ld!o�@&��&�<��Jl��3]��)�3띝��{9�M݂��j'7?�;�\@c�� �|)�������vk�|��%U�'�{�weU1��nI���`By�a�N>�}H�[i�F�i�cʊ�Qr�!=Lxq�Y���Q�	�6�k�>ASt��#�Vx�[�_����rM���1�#�j�D�����$}�&�^zhCH�8G���$ߙp�u��2�鱘�	8�w��5��n��K藪{��5�U���,�y�M�ϫ�ԏH�l1�%n��W3o�G���T���S@�w�9���L���^���p���\ݜ?̎�RWk�lR�v&�1�f��J����t������"7R�}����~�[_ZPx���0��q:'��N�H�ƴ�޾�0����6��=]b��oʼ��T��3LŇ�y� 27���$��B����Df��Y<,�����8���+��,j�qF�DltA@@@DzSQ��ti�.�@Bh��#M�RH�D:(�БZh��-t�'�*~�����ȳ�^�^k���k�XSˍ�8�˚���>>�4�sD�������jp�d�����~��g1���Q�E�''յQږ����1tr�	����tw�P���%['�2=��������������E�:��܃�����%֌Xk���<Op�W� M�K�O��*ś�@nx�#P�G���P�tm�^Ng�0_AJ��#m���c^�zWH0`%��@�%y$�iלP��#`&��h�,CGQ���b�'�9#:��|g����6n%�l�in���ww\&�0K�I1K>Ϡ��3D�eM�������l��_�:b/?+]Rz�^R"�mḩ̌l5���A#˯ uzX�m���C��L��0@z8䬿���J���S��M�Ge�N��G�\�T�EV� !ex���e�#��P/Jf��� J��,<v�����D棤W�?&�'VT��p�hnG�kly�d�"��ɝ��Tk����d��)cQv�	+�!������r�C(M	A�+�r���O�3Y/\Т��a����� ����8�^����ߒ|�Ȼ��sHR�����b[;b��m<NȦc<�WNɾ)���)<��&.�Ȟ����p��� z~n���=���x2J2�@���	^�Q<���١+��T�]��j�q�b�6˫�`\e\������+��}%~����=�<�pƖԑ�P3��B�?����pw���ւ����[����~t�R$g�g�զW�db�⩕�CV;uu��?aQ�d�{�eb�3�5�@@|v�d�҇�y��[%3�o#�N�����#Ȳ�;ճ�?nٚhW�� �2�#v-݉�苛��c@�A�V-^�b)>�;hm�	�U�Q�c՟�B���ik!߱��v��X߫�ͼ�ŷ�8�b=erY��,=�xV�ԣ�p��z�־<���/t/V +۠Q��?������Š���"�\�������=����c^:ۙ1&��l*1휧�	+"��W)��p�c��Z`]��`�dfis��O�q���7��ٌ��|͓6<����ՔJ�����zY��t$�m�?��Y��i���2����#-����\�^ͬ@=���
��� ̞/�5��A��۟-@�tAO{`����(m���K���gS�A՟�F	�����t����Uo��Ip���{5���	� ��,`E�oTֿ����0 F{�L	j���-���BGs'�\��Y���n�_�,�m��㇁�ř�2d�q�M��.�Z�O�jrt����R�US�� ��~��Pzɥ���.D�*�6�+�u�u�F�>��~�ɓ}k��j��Z^�rrPׅ��V7��}��J��h��k!qXd�)s.�%�(�]�늠��,�kg�ɓ�P��t�}B������2�H�*���2$�񈿜plN��\�k�#k�ZD���6:+y��+0��ТЎ^���� 3Xm��6�U�7q��dH`���D��y�徵�_�.��4��(3��:���	�dU:�����g�t�P����i�v>A��2� �(����/�z>�6n�e���!e�����pg�"��ͽ٢@d>��|���˚�L@���A�ϐY%a\�����΃*
�������V�1R���[�҆jn��e��&���i?uwq���W�ϠZ�`:Y�p����z��2���p���l�ԍ̉{�̕��ͳ�#�z�!Ry�{��tc<�:�X���w>C��x��E#��[p�#�#�|u�����~^�����t^���H��,-���څ�;	��֓�e:�h��������0&�/��m�@LY.�K����?�i<�����Aqz�lOy��U�S��l�]�ۑ��%���čg��r�3d�7��}z�NG��Ǎ���F0'p��y��ѻE2����� �]���{�з7�%���\�>�I��v��/o >%<�Taƾ�y�f�)�9��/(���-��kf*�y$_� vI ���(Y~�q-�n���&ɡ��(���jV�?�|�r�kk.x��,�<�oZ�%i�f'�@g�~}q��!�#�GK�:/�H�o�M�o�+�"K��J������C*� ��G�Ј���lkZ�'I]����;�,^�w�hse��E��9gي�G5�����4��x��u�� V�B�z(D5�44k:�Iv� ��ҒX�|��s}�������'�б��7p���ҹ���2�?H0S���x�_�t�a�i��������Ӓ�q���W���~<�$i\C��bh�ju��_H#P�a�ܖ�G1ނ���m��D�3������qW/����/��G��)���ck�*Q�&'��dG�[Iۇ%����N���k����c��g��r�����#w��o6:$�\�h�,!
���2�o�%�ɻ�w��Z�cO,7��b�g(V| i��Ts�ȋʽ4z���ѬUv�jt��'H1�Qk*O)��<�{��|֭�u��ENI�5����f�G-��շ���v�a��Ǵ�u�C�\���;vߟr�+���$��׊5�=��j�����u�@{��.����L���s���	�Ny�B>�����טYF�+�]\TR��� W���\$ae�3L.��"��4�E�#W?<ɞ�Jl4l]�hI4�˝jU7��>[H-Dڢ��;n�|w����:����#n+F��l�D����r�Į�S�؋�h',:8�K�	k����d�J �������髿G�u��T�F�>Kz��ϫ'�/��ˏ���+�;]����|M��x`)[Q[K�~䪦�E!f]
$��SN����E�)G����A��r��ړ	fA��9憉Ձ����B:���kH�ǽ@�C���
� �Zj,f��a�UO_����c|®9�v�h�c����ev�]{���׆1��;�5�u8]3�,�f��y�ێ�K.�oiLI���?����Ox���� �ol����^q��9}�-��|��p�,I����/��K�gQr_�p�1�|���>��|K�iӻ�/�Gފ�l;���Ħ]L&���Zk\'e��ݨ�~bVuGdu+���V��o�*�{�!��M}_ R���n�%!=�U��3@m�2A���e����U�י��j�XW�N�Jl�-9][��K�q�B���,�*���J�K�A���rĽ�H�9���E����I�^鿫�̋N��$LNM
Oy��W������~����oFW��Y� ��o�	�v�5K�Oڊ����Uڌ���u+�/;9v�n�)ޗDw�6���]Rx�<�?�M��}J3��#�I�yOn�_�1ę��>pف�Ұ���<�uϤ�nL>Q̈�ڟXͩ�5�^�s��qQ�M^�qY%�/{�BT]�7W�l̓�)��P��H�����7��y7����O��;t�RixB�j|��K�2V����ń�̣$�.XX��0~��٨ƛn������ﰪW�Kw(i�n�B!�����)u;��^:�n��ą�J�k(�sˉ�)����n�'�e�� ^�ǯ����ڒ�`Y�Ij�Ms�Aō�.�kĴϙz��6s�͵�������<���H�V[*P�z%��L�(�v�V���R�\c�93w�D����u���p'9V5��ۚ��FF0&���dZBgJ�9W�^��b⩄W�ho�ET�"r�QY�':�5�5���4'�S����u �3c)~� ��3�-�eq�8�g���СJ�����6O�Z�FZ|��T�o� �y���� ���#yJ XS$Ie\^Е����� {O�c��J�Ҕ��g ;;�Rӣ56�t�~�fS�+_�+Y[IpsC�k���Ý�u�c��,C%�<|~�J��7����Pu�4�u���/��	<��/��K�6����~gm���/JLw�׾nl�GD������3�#��Rw�Kn<�>���u�D��"��t��{(�*tcZ�D�qQ8~�s��\�Da�S�;*n����ݤK�L���۝њE�Gݴ_�Ƅ�^��~�ǋ�b��4Y����N2ɒ��Ρ5;��n��T
V=5h�e�����,�y��HF��}��}U���@���h�#]�oƶ���VMUEŶ�����yw���������iE�������ʏNH��q�TnM8%���>��z��f|���B�
���?|�F�׆���j#��u�wn El!q"�ϴ|
��{ո0v��{]В�A��H`����fO���{����STP�[��w�-�[�a�Y'���X����6�,�T<4{Y:����o)���>]@ �;O���ۯ`��p�}��X�w�}�Bh�D�|u]Y\;�{��R��']o}z2<���`L�,�粈j4G��^�A 	6ddR=�3�4��u�yb�`qAN���m��]�i�:�N? J9����H�F!�y#	��[��F E(��	�j[���S�����(���y9���<�4z�j{J���;W���s"�ƒ�c� �
��ɚ�}Y� �n���~η��f��k�8�s<�&����?��Ҹ�����Ilg��5nñ���Ľ����g-fW�V@H�Ϋ�/�W����ٛ{,���ZR��{������nvL�e��uwmDU������~�S@��X� �X��zRl�v��9��ݙ,��q�Y��Y�E��4%��ps �s.,�@96L�Y���=~��\���8�� �g�8!�]H�SD�%�4���|S��E�);wїz�]b��;�6H���#fꛦA�V|A6df�~1�����v�V�����C��!&���c����"oZ ��a�E\Ɨ����jS� �G�w�tekq�����m��<죾���e���ۇ�/:�7=��(�<=7�|�p��	�]�9�������'nAGL���[�3�wrތ˲��5�_ѢxD�?n>�/��d�]4@��4��v�/X���%����w�t��!�o��*gL&���a������B�G!8�8a����-�z{��(���˧r��QlJ,�����P��������Nnej0��s�����a�- �-w$�����NE��x�HKI�Q �����Yĥ �D=�N�<ٷU���1x_k�3�ë���
�u򄌹�ྞ@�|O��v����ˑOp|9s�q�O�Kq�<i�h����7y�k"R�@<̋DK���)>`�v{��Y&��#�x-�wR�?�a͋hd��ow�w��.�s2�����<�n?cb��0��b.�t�X럠��}�9���4�*���|͙��f^���/�1��C�`�ke�gwjzc>9~uu�"i�y���>�����l�G�LBȢ\���s
�ԺjKR��`�x]��IխǓt��g(�R�o�= v`�N�� ��m ��P�@�5�������7�;�FD*�V���++�(�q����@T���u�(�(��h&����Q@D�	�Gʙ.n~>2
Y��v��{�UΘ��X��Mt�cM�[Uidq�	��b�Ź�4��yo/����S:e�����z�}%l7�y�z�}�>�.;���2�:���Mʿ���wZ�d_rn���aiڅ=ܾ�qvחB�N{ۗ�y�MOϦ<���H{��C�����y7KC-��d�.w�)�|����-�^��,��������֌�����D�~���@��v�N?�Ԓ�fV����oS�uw~�_����ѡy�/���
~��}�#Ӈ4�d!�tHȓÔ�s/1��G9w�(�e�SG�u'�Mqv��>�feqc��1-|����v�J:<U�*������2��+�h��<�u"�: ����k�إ$48&��	)��\�
ٕ����͞����Q�V���{���������/�s��oC�>$�n�.}�-k��D�oJ�:��ɟ���;kJ2NGqs���V�&��r
��"���B?N����@w�ኦSt�|��aY�Xܺ�JmN}/Ͻ�S���䫙�:�R��Q�z|l1Z�+e��j�;̈~)9��?�#ETz��!TY�
�ހS�j�O �xmE{>V>uFY��n;�L�qnݶ6��]3ܗ1�|��g���4�G�|d\Z�X&�W��%%�dy�ֿx���E������|)���ғ�v)(n�X��Jf����O��M�ۧu�&�;�������w�����H�b��xBNש#ؾ������1�B��j��c;���4�9')�l�T�ň2��ӡHIz��oE(����G�N^�(d(�_��n1�T0o`�_2帰�F�Q��qQ�x<���g9%�6|�U�Ã1( �s��>�%���U|�O�g��]č%.D�Y�Cr)�ɕ�z�`�er���<�5����Msh�79`<��_�л_]�Ȝf�����OM�$���s~o��0� ���{�h�T� �RT��.��
���%^���K9�٦�K�{�{��-�P��r�C'5@3�dOt�ª.u ��%�8����Fֿ��w�|�y.�q��U���G��^T2���<�J���J\�p0\P]*��yKV�-6f\�d�6��0���X`�?�?�P�H�O���	vЈ��_��N�VH�\)�!��8o�rx�O�R�߮�|gہ�rI	�p��՝Oj�Kc������4����^��c�~>A�G_��P��\��A2��>��0P�]���T��>l���+E��Kڦe����6��;��]�'��ȬvO�f����ɹ���y~&O|�g�em(]���"� {���ʺk������*U�am;o�R�?�9���WpW	O����q��n���o�ú��x����s�����KƟ�.���P��(�j���L��^��;�����ގ���s#׺齺Jo:����؆�G1��Cߔ�VD�{��x�l�`�ȳ(��H���W9ӳ��B�1�ծ��
\}�Z������ C�������#�$#_ހ�E��l43�5�Ɛ���L�5�æ׉�U�,�޷� ֒W� j�t+������ p�G��t+�4��ȡ���2�$X��k�Ύ���1�l��ɸ<��� �Ɛb����y{�G�߼���׶*}�چ#�_��P��}���R$'f8*��+���!�R���8�<��x�����yO���l���݆O��fm.�)B��$)C����>���Ջ#���{>Jv1`�xUee��' v������!����	>����W{ޒ��ZQ�����ݻ_����ߗ��h)e��2�!�a������^�h��f�B����W���?Y�#�1&5eX��>/1~Eܚ���Cj��^v��NDke[�bz�j/{h�l2����]��nu=�C��m41�)B��TQD>-�݇w���� IM��ߴ���
H'����L�߅�5us����^G6<!Hi~����m��f5����H��2L���\�1�-�a��gnƅI�����5G7W2L*po��W��ɛ��4�����c�V}Ȳ�
o���-H��"5����R6�0&�;C7� ��{�l���w��B²[��d�$���Jڟ�Z�z��k"�����3{-�~����N[�T��qR�74#�]�;�
5��e��{sj���9^e#B�x�e�]4��*�B�V-����}N��fTx���:E��1�'+9��⌁���¼v-����v(�N��Wx���@`7�MfY��]2K�v�1���^�te���Z9CDDv��cV�n�[������@���7#[�9�2�:OU�42��{�-���c*$EY��A��y���c�^��~^>��������Y�1�2	K������1/ٲ�S����2����;떗�}�I̚�n�ѽ6 �hV��Ҿ]e��q�y��̗Q��9�(|9#�#l,,r�WK�I���;|��e��"�����j
,��| �oTba3�u��KҞ�ظ=5B;�T�� �5�>�#��j��Q�N̠�nEM�ʻ����h�)g�
��o�dV��+�(*bI��W���^� c�͏��$$�+]������ˮ�~�C�u
�F)����E6�'I�z��S�6*^Bx�bl����V���c�FW�2�!���ۙ�2�n���M��v����_�v����G��䭄�jv>]�K3��;��l)2�7���e+���
������p뇶l��w�M�{=�o�N=.iF�Ԉe;Q�v*E��*��ᓗ O�#�4�,�U��2u~�|];[lF��b��!�9~�oV��%x~ebo�Bq����6I'���&1Yp+�F�W��lc��c\r`w��| <m
"�o:Jk�X<TP6>�����s�;�W�,w�������}��������kP����ԛI]M�4��Z�O}����A�8���澥d���`2W��Ȯ�^jŀm����3[$�	�t ��v���/�6Ñ��:vɻ���{d��ҏ�^�-$t%JED"TQ�-�g?8�9��"{t@��Mh��,�ڮ�ݚ�6R����5�����9�TZ4�\���p�e�2����N2�w�<�4�o��7�;�b�.��*σ�c�	�����~���ÀC����l�Ҋ��#�2�A�l��X���d���J%��k�痏�>�A��={��ۛ+:Q0�����>[	\iY�2�5g(���cS�� R�0�x1��t�-��栕%��	�	�{�BJ�`F��y��b�����|�^Nɻ�a���!���i�7��7�$#��K�����MQ]{�;�^�H�G�)��D�������	�����C^��	�p�{��N .�5i��#"v�Yt�
k���L����.v�U���w��{��Fj��� ��(6��M0�X�W#��hWg��Q�H3.�5x�Z��W�V�ri��/�<t��/<���>�ɚ	��0ٳ�7����BE�L�I�N(�ǘV���HꞳ�R�ܤ�z\iD�]"�W�1mPdn-�W��m��?�NF%p^9&�mX����R�I�t� ��:�hJ�VԘ�'ܩ�Kg"��Z}xv�ɴ�eC��;u ��,�y�s��"׵>�b�s} �9�������`|臯��3�]D��#��rȸ���T���}�hEfs��4�ǖ���{�j��kB�L�Y4�'�?\?�X��UW�a/�7�ks��2T�ݯw�ӂ�m��cK���8��$�ܝ��O�$
?��|�j~�#�/h^�����2 �@�*����_����YMw�׍��K8{*p��\�����`�����@��������c����^��E�^��b'^"�S!�0(9�Us1���� ��I�krk��z���-^��k�᛽�1�ad*���:\���� �q�ܹ����}G�}�+�/�i������Odk1�	4w�����Wi"X|�ݵj�x�yh�F�|ߨW�|fh#
_��_R�gd��MnaVhY'����#f��J��}4�x��TD�&�^۬��@)y�Zs���t�xw�x��n�#M�����:�d��4>�����]�x�>�7֒��)��J�B���}o�h�V�X!k+�/���CT끡��K֡�K-;���nx;��1����|˽�c�ɜ�P���X��JY���J�&HJ"G����jоu������W=�����h�]d�{���֤Ny=���F������2�X��&��]I�t��8U�J/�^fm};���(lzS�E)Tܺ�8��U��DO�H�*�c�{��l�PF�C���Q�I�MY�s�lV�%�L E��(ĕ>�f�6�8�jｊ��A�������̆H������bH��p�˓pM�̧�X�¶�s��|%�|�Ȝusc��@]a�#���w�RE�嶽i�|�1e��eA���d��NrĄb4D�$�8��Yl4�qd��^n��0���Z�j4փr���so����^����^�	���}L�>�+�,&��Z#ӑ�o�/g�!J:GP2�V��C��l�ƕMYs/_�%'�X%��EV �Hd|���UR8�	�=}�\!�!y�M��أ��n�N��/nƧ���.�(ź�r�h�]L�xSSP�h]�(f *2聽���@�p;�w���ķ�&�Z�C�m^�\��D��Ț��/��J����OOrw-P���e�!���M�Y��"sr�>";ԥ:�ϐ_'fG��N�[�rY����\���e^*�����i�nn*&C�.E֬U��ͫ�Vt^���Y�:Vbߍ��J�(+�[�!�?C��뺏�H�E4�eW;ʖsŅ�7��v�,^}w.E�����W��h.�u���5��Vr����}Q�A���212���̙�M#s�&�q���d�:��f�W��S�l���`�ė��sk��#|��麋�1'MT(xش�_���A�廲�F�f����>O�^�W_����o������N�Ds(Ją�">Ď�[tT��e���'���u/	��OӐ��h�^�,���n_��lޫ}���4��e}ޝ��V�$&z�c�S�K�-6��bv!l��p:�^�ǹ�2�~�j|��^M�ػ��}��D�8���v]�\�E謊a&�1l�ˬ��4��~�?�k��|���Y#"wi�I���/˖� 2���Gѕe�R?�Yx�D��K��2��(%EsB����f��]�ǫ�"_��R�����:7we)r��ً��vB���׮Wc ��h�[v;��e��oS%�N���R�Aη����8:��r���j�m���=���,N	��ފ<��47
�hʼ>��"����T��&�p�,�f��y������De��\gu�K/YIn��׽_�E�� @w$O�^QW���2�@��1F3�􃓟fd�ܹ�P�
�hٟ��v�������+%�Q΢���d�;�x-��t�w�TrE�[A���N���F��E�`{_ҹ�_&���$(�n�n~�XL܄xȍ���w�M�n-}Ѫ^؉��[��U�=�����_���J�l @}���b#� s��k�7�����x��Ce�w껇˦v=wH������E�cϪ;���������]owP�W�,5W��|t��i��#8iT.s9�}�{x�u�&�v���l���}��7��GPV�zc������p$�5��[����vF���[ʆ�gj2u���U���-.,I��x�����c��|��br!�ËoY!5v�c��p�w6h��r�Z���49K���:���p�w Svy��-���2��� �{���"|�zRa��*����G��&rl���S����d4��.�>dd�H�"��)�C��H_	�l)]���ś�1%�VHl�7��&��j�|��k�^��>O����ɇ#�.�Q�;d�H���[]������XvL���xjc�H2���K��.K���*���Eσ���=����U���d���v3f�I�}V^���׹"�,�y���a��o�0����u��[��L��%qG���wj_y'� mc�޿DrX���m���,��2��Nn@�	Q�p�R�_E92*���.{53j"�ۓ���d�lʗ
^Vz<��R�<3�/����!�]���:��ľ!b��D)k��P��nw5�4,�#d���
�����g.YU=���vu:��0�	u J���� me�:�ZI���+a	�F���\���ߵf�����Y/��f�5��D��Z�'��ӥ��o�DJ����^�YeM�攗%>{��<fN�'gTV��1\El}�$i626��^uԪ(힔�$XDNn�#}����I���
�_f�ɽ��b�C�A�&�h��[�;F�r�����f�t��B�wj�M����	(�M�!�dYT��dZ$=!���ӻ�C65T���֥�0���}���lb�|�_��;K�r�Q땦�s��� ��o�1`�j����ڌ��2|�ܞb��K$����aG��ꊳYn��R_�)zm1��b�Z�����d*D���t�>�������Ϻɍ����#IN5G����2��5".5�0�./b����D%�vX�N(76���U�7-��뺲Gϭ��y���{$I�:��������V�ƍzF�9vǳ����9c� Z���NYrb)��'�¶%����w��/c�ݠ���G�%CM%o N�;"���GH�[C���A<Z܌��|M�����2����S���Tr�������7��sQIѐ��\=K%W��Z����K߰�@]+6�o.2�']h�%9w]ZJ��4���&6�X�%ڧ�V�/������2��@�]VF���k3+������˨�PA�ʛ\"�U��
�]��nfE�y�i�uC��l��뤫��]�����e7�&��r��[痲��>�y���D�K���NX_�&Ķ���v&�׆J�s�hxw��]\CI{�|gq�� �������V��i�b�_�bܪ�_�;A���4���J�r~�>��mW���c;.�.N����c��0���+�Q�z�_��U�P@>�j'� �ti4�r���e�p�R$��=���m��'��8"�w(���|�}����ʣ��G�o%��7�$4?�?���S��U�iV���MQq�'24��y�s:[æ�\��d�1�c-�T^~�N�k�	 "��g���}F���~ۅF�'�sױ��s$d�sy����̗��٢7���� �k����6�.j�ܓ+�H�)C�	D;x��4���p��"[�x��W�5�;���Q��T�;h;�~R놕�&$%�=+�23���N��]���\��.F�胚VĉD��v�A2����%5��ؚ�'� \��v�\�����F���S���<l����Hݍ_��d")@�Mę��`�T���Oڸ����{++�i���NFW�5��r��
�*�&$\Ue��k8w��%��)cW>@d<r��I�l%}��M��Z�R�8�a��
q)B�@�r�:I�����J}s|�`F����EXa��[�Ee	�'2<�.)�5������	V=�<��3�W�
	!o�>I�`�J皋tm��cl1�1v��Rc_�4�)\+4�Uhz)
��%��[���(�ATd���MF��I`l݊A���*>���d�b����Ӏ��`��(�.����P��U9���@m��)˟�|���S�V����@��{a�K���e XC���Y�x�ڨ���.���{��L?���3�z.d�)`� g����ZI�P���G��`� �-k��K9��WJ!&��L��yb,�ᅬW#2�^�:�J��LW��1*8&0GÒ�ͦS"A��f�=x�WD��*==[���{/��T(Q���wˏ�����K��ԡ���@�����:U��r?�����@�J�<�0��h{gnd��j삒���u���������xۉ�v��ɭ������O�1N�tC*����Q��������y>DP8IU�����pO"�@ї4�g�Vy{Z���8�'A��D@�Ce�^�S�	���}ή�H$t��-�GE����?���W�'/��Kbm�╩+7?hx�hU%N�V�)���#`���:�;^}��B��ϧ:�+���[ؘ��C��KXb5dNMvS'>�2������q����J�����{F'7���QK{�M.��Y��1"�>�e��s�h�\�����_�A��ӧ�kd���Y*,�Ҧ�ɌN��_V�j��?��>��y��2o'*�41>o�_\�@<c�wU����ڔ�߾/R����ԕ�l7	`(��	͗,����%Ēu�ߺ����|�t�+Z���d؄J&���ΫIl���*f�}`�+���̬xç��<.��L�(�\�����F�F/���w��˄��2�a���fe�|�)����Sj7�y\���`e���Y@�N�����/iΚ�2��6�$�bΊ�*2�C7L���y@7��,��p۰� ��@P;��I�o	ղ;a*�` �..��<�0&|�e�-Fk�$z����R\�a.��U�?&Ӡ]���*�����G�c��U�N7� �/�:6R"
T匈Y�^����W����>�N��*�I{�ʇ���в��� y�"k'%k�8�R�����6,�MR�5�g��i	��j	��7NU�<�Y �����5�U�Z��=�ֹ��/A�`ݾ=)�&O�ơ'����u@��0���SA��<$��K���8���� ��1��ML�_��#+j}jz(c�"�@�+��ǯ���%)��k�PA���7�S��[1��t=�E�:P�_~��T���:3�QjIŌ��D02�)�Q#�3j��ٚ¥��|���A�E:�9���N*;=���>$������ �u!��*�?&��h��M�dA��st�=QpKX��h�7@K���M��`��,���x�ύ\J�j��J��Q	 g���y/�r�n1à4G ��4(�J�!�:F*�$�^�g��cVė�eۛ-?e�J����\	�<����������+��1�JIe�j�σ~�rIn�$��K�J�PKv�Aq��VD�c��u"����W�1�G�����5!�nWx֖6#F~410A J3�7x�R&�HFG4�(��b���w��}��[̈�f�t)��g��(G��s$y�Dw�� Ee���(;�QB6C��VL�~�[�رf	\���Ɂ��b �H��8��o�"����&�ߤ���*72~)����Ç
�Hb��z�1�ʡ�b&�wJ�S"0�?�V��i����XM����\aN�+���+w�V��J�݃��8#_�͊��V��_��	b�/:��bB�6�s�1�<c(��O�!p�HPm1�w��oZ���"7i..�م���}z��ݣ{�����i\�c�"��|�=vhj:�z���al��¼#���yF^��o��|;��1�h��'��=��Z�'���|��ۄ�XFJ�+g,��@�P������PX�+��T���b��mݖe�m�w�F���jWÂRZ����W�"���SϞ��/��w��ߜĳ����#-,�������l��������_Ϸw���|�_��O��� �_N����K���_�}�9����?���} A����Ƶ.Ϭu�)氺+���z�ؽ�\���\�����K��C������T��n�ogg�́��[���hRy�m�$O��A�Z:��W�_�FRfT���"�c�'0� ��G
���(e뱉���7�G;�%y.|@��w{A݋S��T�["ؐ�گY��h�:,��:�H3��OىB�?�,��0���>��˝5����?�� ��r̀z�62�a�%=U;�W��
HL\i@u モ��52������)��������Z�/�ٱ��̋�b��5�+-6G�
5�����mUv�iU�j���������ӷ~X�y � �8���+̮�R��6��buu�#�w'2�����,Q�_u+2Kʹ)�������e���-���mDҥU�2y�Ld�0!���V	Q��c���A2Q�N��֠�6X5]�Jx�M���3i� �{��F����}v�aoq�BVSp����BHe��`r�����	/��ێoJ��U: ��;:R�u��������u�eyx�a�0�+R�T'z��S��ɧ@����9>`>��(_Q��a��Q>/vſ�N;�R�7cT�^�����1�s�)\�� Ȥ]��W�t7w���@�h��B��q�VG���Q����ny@-�g�����)Z�U������	7¶b�j����7�W5ͩȠ�����������P&.��=��V�M�]��Udh�y&N���w�?N6
�� ��.Cm�H���� ����f��3�I:8��������T�)���.pN};_�#�'�hM�Y�&��[;��潌����P��4]W2�D�:�R�������I���X��Oo�(J���y�륂>��K�����!vI�jyfgק�m�g�/�N[��� *\�/��ч��nY��� ��*�v�*��D�%�=E�^l�x�qB�p�%KL%��_|VW���(9Ww��:�G�РO��g��3�T�'���3�RHj����'�\�
�nZQ�N��]R;C��/��Q�+|/i�q�|Iw
ņA���������.vVsrp���X *S^V���������X��
�8O}OL�=��]M	s�D	��M���C�#c�뻀z�L�!�m?��9�)�n�{���ي���0d���^��m�����M�jxB�y,�nH:6VJ���]r��&»��k^���6Q���b �O����Q�\�sq\��P��Y����Z-B��v��P�d/���V..���fwJ���Q��G��ռ�X�(�_�#iQ׶e����7E���k$~���!$f��h�d�x��>���F:� �l7	�Y�0�6��Y771�0\�Lmq��������7��i^���:�슢+�x��s>f2@�z���r���3�*Nl���t]�VǶJO3WQ�(�7^�Y.b#C��^�ȕ�52��ɒ`�M�W�4^?AU�iw>�(\��q�ҡ=HjZp5�|Ѿw��2����w5�h��\��|�p�ms�f ȝ�D$�l�D�������)H��CpW���~\i�9ŗm]Į�5�����a�N�#�ty��?����v�h��=�d�����+Л
|%����~��~m���\��W��N��O���Α|}H�����
��f�z������Q�Φ��GTn� �� �J ��Oz(��@I-NLp:&I�:LB ��H��E�7M���IL�����W�3YG�~���#~�f�~�^�,��}�c A�����}���E�$6�'�D4��1x5m�726iu=�}s��DA	h����C1c��ws^/g�:��@��W<�����G�n��鏔Ñ����A��\�oR�*� J[K�v8d��K]��V���+٦~OkgLd�ifXh:��]W�D��bOK���P���a���=M��cf<�\���L�>�����
0�?b�ii���a�WBs{6I��/G�z���)hE��p�&�P����VE�}{ۅH�ײF1�dɾ�������Zv�Q�mP�gƾ3!�����|��?�t'����k���u߯{7t��@�smT��s�Ǿ�7ý��z��Q�xz�7C�C�Ǚ�*�9��j���Ů�t�����k��������XIK���쫍�"���*�\۞-s]����N+��#E��}R�}��^!�4A��~��2�	��K��"��MZ����gFRN�o�j}2��&_?�Bja���E5�G6�驶�Ȃ(� ,b�gB�FA��/돓Hn��`�넷p�-~�O�$�&���K4��#�K�B��2r���LЀ����?I�\�V�#ɵFw0�lS}'P=�.#�����p;��Ј0�"��h�����b��3�)�Y#�Tw~�Q#�� �x�}��-��"gF�
����{�^�Iq]��(Vi���O���4�b\d3I�h�/���ۓ��O�;�# O#珄�V�o�.е����J;F+�3AKE���u0B9��,��URRY�A��/��t[q�a,p9�H��啕�U7s>�<S�����G�����4�}j}���$�a^�ȏ��4+O�Vt-V��*�x�',�%	����J�hNr�5����\pnL����5G1�3x�'�Pl�O'.���-�ϜG� ����wR��PR����5'Sӝ]1�܇'.ԏ�i�XR8ACM(#�H�)���Ǉ�	���*�(����?qW̟z�<m0�"�i������p?|X'�;�3�[�'%ʝ�Ӻ�}�s��b��H?�ւ�E�ԙϪ	[��0M�nH�O �h棒�ְn,< 'R�vC��d��q�J���	���-��c��vK�o>�@�{����VL��L]����z�����ia�<���/�J�c)8�=��1"�ѫ��c��1�F�߭�}�[�������p-�6�������!�H�i�W�am����h�����yJ��E��do��í����V���+1]��=����]E���'��um�;κ���ɱ!pK���U��0�z΀�X�\��PՔ�T���i4�7�ۗ��2ϥ�Ҝ�����p$�35�@��,��e���r�Y�Q��Ћ4�a�a�5����0��LU՚ͷJO\��L��3e�%�^�>�׀���;p�@�"�H�����Ko�l��	H!mjE����v���DT�c:|T�*4���I[/���g���`.@�?��MHmX��x8Q�6�9�hk�"�=�����e3dW�0.��|/Y��w^�PѣzCI.ح��짐!x!n�ЏV43Ӫ���1N2nw��۳�]�7�)��G�35.L-��'FN�("��s���M�-��V����5#뫜��-ǲ�;�u�7�a�5Bj.�#��R�cbzn9&q�Ep��}(��D�`�nw�6���e�1� n��������L�?��T�Q�ԯus���昖��4��đYE؟5�b�����6ұ����.�ẾA8�Uᐚp$��n��H�ظ���O������YR�b���s�dDƻ6�(/~
n^�)���RAp����U���Sdd#O���� �e�:s�$��c�f���U�j�Q1�����F�&���vզ�|���D�3���u#��vzNQ�-�ٍu��=��6���7Z��c-��dk�)���f�?���b�Q�&[���-١� � H�7�֒��(����u�s�@�g�k�wĎ�M��~9�暴z�76���&ǚ�襆�);���
>,�����s-ĮdF� ��I�U����b>W�М=���J�c��m�XZ�_��M�J�ʩ��M��;�"��3�m�OT)��E�K����?�wYJj6!����I���a�Q��G�
ԈteW����0��W�WT�5�������A��E�"�*1��T�T���A0������t����xݒ�ӞՄ�3Xa;�8H[��nZW�؈;d��D��:6w�;��ݳ)�ӛ�&�+�P��1�a-}l�drӆ߹X�2��1�"��彡���k�w�a����H�;N�H�J9�t�����T���!yF	�)��Ԧ�Nx���zm�g3�6��o��Lu�(����m0��7~�DL�l�P9$p</�۩��Y���l:0e���8��R+��t2r�q1�A��`�������k���\��f���v�;S���
�2���@��eR��-�4J��KCE�G�W�r�8�V)}����p�lCs�h��>����F�*��	luh'�x�`'�W�v!y��۷���L�U�@`�d�����*B�i6��O V�b<��F�?�-�>M�눌�9�b�	�2�,�tD�E.�Q�z�f��c]�{kkt���[�=.܄��8�o��������k����np�_�s�N�I���o�]i!��|�H΍&�H}�J�3&�s�� �ܟVa��#O��U�3�#=)������6w�+b�"�!C�բz�R��:���)z�����k޼\�l�M��ֿ_��eN���&|���l���?�"O��EeL�&mb��!G3˾�G���:'r�������r���y%�
�uw)���+/����b�ޚ�`���ղ����s��b��jD���je=�»��"1�����	+m�.���yQߨ��\�t0x6.]�����/����
�μL�t�s0��S��Ö%+EԜ(�?����ձ�k:�;��v`��mg�x.���������"2�!���'��0�~��g�!e{� �l����m\Fqs���X�>Y/+0��t�ct<���� ���N���[����
��3E^�]]9KmW��a���N�r[�5!M�O���z�Tbnkұ�N������[6�=�NFf�U�{J�v���"��Et��z�рl�[õN�Y���U���N̚���C��q�k6��<�}��2�=f�.�۲0?eL�]�@��i܇5*ح�&?����Q��6�tWLd�V��Z��z���>��"����6��E��:��bV)�D��h$;Q��\$�Q%ρ���I�j��Ww��M�y�%rwV�W����F�x4��k�,�M�t������=
��l�����?�~�>�8\Z�O?��#H���ݠ���@�K`c�[t�
���4-�ǎ���KWK��
�uA�¶��]��¯9z�y䐗Q�>EESo�70%�8X�T�[6١
8bG�r������ig{�����>K#���3v��)D5�c� )R!��յ*��Y��KJ��{G=T�V{�9� ֫Jd���u�̧�+-��;�N�p:Ƴ�5���/�{��/h�ↅqCV��X{l�k�"@�"����ƱEb�UU ��\���-H�cq��2��\���*C���>���F2DP<�,w㏕5ew�qc���T��j��f� ��mG����Wa�1P�Dİe�2��h-t�
D?醉�GL��]J���~��ҶC���>�H�[��G5h���8t�|q��o�m��tu�%T��f�f՟j��PHzٟ���mZ����h�^���O%t��\M�6�zGD9�{2�����ɧ�_o����^�~��"-�: N��?(��4���$��Z���u�6 �A�bxW�r�P��<$�b,W��A x�aG�V�`�������Ůڏkq����(0�v�E̍�н�p��e]��ďGV������\<X"�V|�! ���}���
d�ս-�Ñ�� �[�Q�`
��nbU!B��	IͿɓr)�V�5�2l	��?ަq��|>���zb��������p�Q;���5#�Y��ǹW�������Î���3ck��>��
z��ހ'k�S�j�yy�znk���M����lu�)P�&S^ZJ���[*>~2>/�QaRՒx�yC��o��h��^����`�[Y�XU��ts������!�hL�l	����@%)M��˯J��h^���w!���6��J��'�ax\P+��@wk�\[�=Y�?~�%*�|�̞�Ș0��2*�۪x���Y�N2a���Y�d#�#�~*	�>�6N�}f�o�@��9���k�M@�k�Yάel������k��4���U�]�M��3�\���ǂV9���̑�zSZkl
qfo�jU�e���,�/�B?$
�߸��C_v��KD���D��S���(�ù@mߝS}-�ma ���ho	DZ���>���0�Ր���3 z�1����d"�~�/�ڊ}�Wc�"CPڨ]��>��q=���Y���nA��yl!ߚ�k���}O�ɢ�c� ��v^Lٳ�7�e��ʾ��k���I��T}����je���P�P=�J��w@᷋�5Fpj��گZ֖Z�����q��Nn�jR��(R3K����8N��"�ntD-,Qb��6�ʷ�8�X�^�:��!-�';�����0�)�n2I���|�@EwN�!�co�ڝ�T,���mTW}B�� |�&Y/�+�z�֤�T���Rlwg�̶��W)Z;Y�nT�͌�;�!8�9��Y=�='��%'�qI^�X�So�k��Պ�FB��K�o���%����f�r݋��D��̼�����	d��
����R%_z
)�{�$9���{K�)�ɹ�8�����e�L �k%�������`����S/�өZ����uH��Knbc�"�7������t���ѐ��Nun���g�˽�Ah���^�by���5���19���`ߚ����Y�DD�Jb&k�U�B���8~�Vh��2d8OZ[�����?<a���x���:s�R�D��'�uN#�k	����?����b]N�­|R��������{��m��d�^C�05MOW�iI4�a)OC�\���:����w�Y�8a���u����}S�?�|X�H�(I4�}���'4��re��]���pV�ԣwԃPp�a�B���CUl�w\�������F&anT�]��4(AU�Ȣط��A�(N��lrZ�٬�.5�FD��S��f��2`끱P�oŝ�m�}+xi3͞_3k�2��.�>Y���Kŕ:�~�W���3	���a�ԧ�
�*k�r���WR���,\'{}�ϗpϴ����/j�^v��?|׫5A>n�KU�B���o,tj/��;���=
oV9�mޓ\����kt-S���P�k���s�Cg\9��Q�j�nl	-�춲BI�����W!�k�-�����Yp[�Q8���xU/�����͞
�l"��ݮL�D��,�X%��#���B�����g<��g�ጝV���M�)Tcn��Xy�^�-*X���dծ��]��^ط��� t`O���k)�5��B�5��M����ɵ�����7���bT��S���� `��J0]�P�P0�����P��/u��OOVu.�{��j��r��,F���\��6!!*��܎N�����$�{\��ب��<�I߿���'���|�kѯ"����q��:.����=�o=�]FF�nR��e`1,�y�s> �.��sb?l�tn5TP�[�^�䉃W��S:�����J�+4�o���{�&Y;���  ��k��s{��M�����_�y=�t��*�Q�>8w�w�QI��\ց(��@��y�R�z�MJ3���?��%)k�^^�U�$�i���l�A�	�r�� e���nC��|qX|&y�C=̅q|��3	�Km�E2�B��5W������I�͡@6�f�B��SX��}�QT�s�#��v±�¡�q���a�	�.�%]J�u�>�ì@m�_ÿ&+&Bͱ���'��[���
�Z�Z9�)����
7�*r�׼TŶP֠�7�*���I#ب%:����pm��ހJ�}N���U�.��u�^;�o��K�,~-��F��~�S��QgqN7\M΅g0g��������K�F�ل��%=[GA�b��_��15�R���/	���ڗ�"P�1�����@ �ș���%L��M�Sy��br<#5U��7E<^�n}ۀ�(�[#g�:�J_u#�p%xj:�"��.�"3��UL�B@׊Ӻ8U���tk>����nb/�5��|zKF�x;9�T���r�H!l,������e��4�/����o3�@0HK�CK���.X?]5`���l&��BB��(���������9٭\��,ӭb�_���%|ZA�I�ĶrR͖7s��Eҁ7`����^F3�ŏ�:�{4?��L"����L��Ǵe�|l;LB!"�"�>,�w� 2F�l��I�3�B�E�7P��n�7-v��!����];����p� ��pesG"�qv��)Q�����h�U
�!F΃M'�Z���)�Y�{!���C�>�����W�qh���Fڀ���=�[*�D����o�Z�`���c>�ȱ(g�܁_]�8��9r:�XU�zw�d�3�ݢ��6��~dDP!qش� D�q�K���#q��������^��-v�8B �6kPt�xT��T����N�
�7][�(�g�U/<h�5Ƭ��;�׬"�G�� �=�M��������I�iO���u�]��>����"���#M�Ix�|6�v��@A$����
y]Ie���^��I�C�j�˭ŏ���"Z{�ް'��һvΓwn��ka<�t���t�=�?��m���7h%�B��D��3R�Z!#v�nS���U:}X����y�{5>K!�U�)�����yYI˳,Q<2:|�	��0����w8Υ�/��.b����Y 3}�A���C�`����t�����S��W~�����;��_��r�87�#(rFxj��ĺqE3և�B�wʘm0������O:��:ǖ����z2O)E��N�� ��r?�;����n�fT��l*{�w�$�*�GSV=֦/d~t�A�E��T�q U���Q��Wϒ������>L��f�b:���(���y��g^����'���T���i����oN96�
OPR��
���b�>E��>z0�g�����S�|(B��տT�?3��s_���>��Y���O��?��900��[Leש���� �����#X�J����Ϊ�4��1�5�q����բ�����}z@v��u����@M����KC�=�����Y��J����`��It��)�sCzNvQ�*2}�scttT�>M��p��j뚤�TU�ߕ�F����o
/���V�N�4'������ȵ����U�P�;���'x�E�OO���IX/�}d�-q.�hBB����|���-t+2�ĭ�i.�=�L�!�# ��Q-�<�ޏ��(q�0(�γ�th��*�ʫ�ST崚�6���M�Hb��'�'��q�g!:�y�8+�g,: +`&�r�Y�d'f2�O�Sf�"ѳyZ��� t��@�'��d����RQlv�S����-���7-�++Q*S(�?��n��v�	��Ýo��*$(֯��?Z�Փ�5KZh�o���k�@	��i���~���6g_��3�8�}����×��f��8�a�,b[�'m]<�M�w����a-�%`z���0,\��;6���n�梻��YS}
{�t���NAי_}Ē�j������B�^�}&�b)�G4}V}W�6(� l1c/��{����X�מHP:��M�A}�����{��@RX&��B�~2�-�Ǥ쐒f�y��Q(DZ���o�z��5K�)^��\_�uߤ�sA��v��#�| R���w%XD� d������D�:s��?=��=��N��/w��O�39�9�+�l`v���p��1e[��h��"��@#��Z�ow/*�G� �^�0KKE���w��ޮ�ٿ���yO��V�Ǌ����/Ҍ�L*:7��{�O�8�Z�nR�������.Vb�o�pm�UU�b�sd*܂�ސk�/i�2��e
}&���I���y�u�zY�VB��������f-�6V��Hq�!��X�����p�N�Ƚ��cP��+�0��&E:��(�~��ƍ�Z�E6x,o��{�H�cI}^�Lx�̿��"��,���la6���"�c��㝃ݞb�i�!(x� �N�69w��a��!�z����8w�k�dj�D�걗Ì�-�h��?R11EeWX(�5n�^;���sfR 0��ؘ".N�Ȉ\���[�u��@���xv��'�[��&�u�IK0b  <���X�蚘�u8�{�,�:s�0v����v^�a�
��h�4�}� �,�Y���"Z�"Z�7��Ӹ��ru<?��uX+��_�m���ԟ{�
׍ c#{�ގ���z����:`��+���*D5EwKqXQ9���\�Q�pWr�Y{Όg���F#�����|����9y�j�X���D3m�1���";�U�J0ݸ���*G���&,���x'y��V�`����_���S�q��e���F��Z����m��:���#�q�C�F���}Z_f���:��B��xw��)c�'��%��+!�<:%��񹡊�lW�4Q��U�k+u�Pמ�z�X.[�j{�vv��"�&-\��]q�`���]w9;�^�?���h�]�W���oc�kV���}���T]-"�dQ��8y�$+�1�/S�g�����S`�je�<d���G������QGu�Ƃ\~9�}r��"����PW�1wVE]��*���� ���x�1����S}�+�l�wC!c�p���s%�`����JY}�*����D4r|�a}4]�X����!��}�)���ȸ�<''��5�u��m-@��!%γ*�B$�Y�a��nH9э��p�Ϗ��gf.�����@넅�Zj��Y��D��t����b��J�̽:�����s�㯛Πq��"�q_����$Y+=w�~�Ϩ@r��{�U=�����PO����K��U�����i,�@��86�c��hMW�y�-O��J��d�L+��%�_ސ�n�x>�mjJqǘ/�7��ݮ؏j*Ї��{�'{;X�5���q�m�K놸I���ߺ�2��5<���_�L�k>m�,�m��j��	|2Ρ����\�s�^J�L��0*{�S�ޝ������0����Iá�s��>g�e�����c+������$�[�H��p�h�P8Uh|��M޿�/_�?@��_"�� ����~�ڵ��u���4>��X��)�7��2���Y
>L�u@�^���|ƹis0��81�a�;xM�g���D��oV�@�Z��O�k�dE��Z����%���?�d������0sDG�^]�t�͐h����fɵ� É�A0J��ri{������'����K2��lې��T�=(e� ��o6�Us��[��j\�� �:!Z��T�2���=%�"�ٯ��/L7A Ђ���|���nq�lѐj�v@��Z���Za(��s�RZ�gޤ�R}�A=�M�^�<cd�-��Y�\�7��{{�
;<���������u} ���Kz]7Hl��-U��z1h������&1w�5�*t^R�R��;8�6���8O]$�ʖ���R,�B����э�o��ص�L٫V����o�o����H�V
;�B�D���V��B�#�r�=;��G�C�ٝ���	���L�{7���b3�2����Y~�?ud�H[�Pk��oU����������npU㪔���O�_������Z�\_�Hy/�m�'�S���w[�~��*NMd���f�'}�;`=��i�O��D���3; ��]�>��@�{.br������Dް�*�:��%~C�U�a�U�'h����&}���X0K�b���	/C�a�Z�ԑ����!�B�K����6Y�n�5�7�h��J{k�D��p0e�?���vYA�%���ӎs����+J�4�"�/4��@�2*:��#�6=���I�WI`�}��g3x!�V���Pb(��?��8����42+߃�`MR�� �kNw�,݄��ZHzoÒ��VGy?�ey�7(�=�.r���W�OIe���J㧐�+��{ m�w�v�n��Q�V
�S��*ٖ������^3(���(](�]�;�������3��N\EU)���gW�����g��=DV{*���d����zI�e�6���,�4��e Tֹ��qn���G�˛��*��*�|ͻ�3y�4*;�tq��Z�.�-�Ѝ�r1�z_3��R#bow�e8;�~b�H{}"���zx�}frn��d�9��sϬ��Z�(Vd�B��(��a��*7���El�5��k���#��M�Z�	�G<�kf{&q"��7O�(�WO_���FZr.2�?�$+����yM$5R|�Φ.�:�TP�[Ũ/�F���
��~v�I���
� � &�+_n���:�2�1Z<�*�h�J��c>Dd�~9�~�Hge):޻Ĉ1(,۬�<u�P�D򼏥|��ִ�K���E9I9_�o]���-���c^�<����L%��l}ڀ�\*�;X��<3D�#t�]^C��6E� ݤ�b�ö^P�PE?�D��GZ�b\�^����9��7P�暨K�9������,���.��β��9���̓�z�]�ݽ�m��Uf�Y��4��̞��z�|d��/a���=pgяiKڱ���Iz4��@fJ;cV}�(C�3��P*Wun+��1�xL�L����2.��y�(?��g�HK�~�Y
Fo��� ����J���>2`���_����߀�S�}�J���B�7��Ѓ%�Ui���:L�A͉���=�ߌaW6�8�E�3���&mV_(���
��}bL�`sw��.ם��89G��k��D� ��ð�����;d�9�lo_����l�b6�s��x}�J欠�������� �j��'�Ѩ�������o_6�PA�0�+Ч�!æ��=D�w���'S�;���䜐z��R��	� ��Xt���7�U�L�ޔZP�XS�x�:�D��Io9�뮼��
�^���3Vzi��Mb��@b�e��2�;�Kׂ<�۾^�6wtn=6~!�E�m���Rx��`�l�v��<�@������c�xh����6 �V��8��c ~E����;��7<�]`�;Ys:�_��+.-Rr�������S���#r��R�W��4�����3	MH��=[;}��4#i�,Y _:��7��;�;�Z�U_�^'1�G%��?�Cк�>|�e�Ξ=�n�=��	ZuR!�7�>��h��ϊ� �_��QSW"2��߫E�Ջ������h��X�	ԙ�*@}�
��ߣ���I�&�=W"��s�����VD�B���xҪ]d�5�n�n�<-90�T���$�E�g�@�L6zUۡ���.nrw�jd?���'�~�<����r��Z�n��)i����q��}7�=vˉ�� ����2��(�QK&��t���G��̈́n_G���i ��"�f-!s�o"z�(�f��*�ؗ�L����e����w�h�<{nwݬa��R�B����B�P��zIc�:.�"�U�N�{�j1�:��s��g���)(۩�ȋ}^�+��0�h�e�!�Ȉ]���;�qeJ0t��k g���>"F�1�n8�s>@X-�3�*��?F�^�S���g|y�@�JjT����WZ�4�d ����'�tgy�B�P�F�3�&�����O�|�]|b�
{�^��] ���
��^I?>a�!S+(��ߗ�W�����Ql�:U�1����A{l��/ǿ{,�/ȅ��8s2�6���8<O��&��������Un�W��:%�G���NB	�L�E�j�4`�Yd�C}Rrs�J;��mBB���*еa����_� uE�9Bʭ�m;�Ĩ�*v��%�{���y����q�Y��D~f����}���!O"�O2#@�Ű�7]���P��Lg�:�Ӟ.����-翹O�5�����P��C�����]S5��.O������i<R��'�v���RuD~�2@�h&��+����[6۸����.�	+�BL��{����P�K�4��3�0�o~2Jn�޲nӿ^�^5�;E�㍛��!��z�}��<�z�����E>z�X�3�Rw�[V����P� ł�����/6?�P\�;�}..�HH�,�/&5m;�$X�W�={yib�i��}|�{%veH��]�ݲ2nu�V}ƶC��;�S5j�,2 PƮ
kѸ`ٕ�d@�?{�C��U��n���*��K'�8]/�#�����68�#�����{[9`���뛇D*BF�m*�0#A}��Ȕ�6�|݇��gV�@�����h�U�@Q��U��E��SF�
�}�[�\�����b���H��+k��C�ތ��,�٧A�&M)U�BO%�N���`��y�g���Hϖr�C���/��Z?氪9F�<ԜOr�(�W3�� �M�ǚ\���6��)��N�w_�gv���N4��5��W��_�CE|Z�}�'�U��G���2U�K����qn�����P����!�.�ڊ ��ݮ�J8;��A��5S궻���#,� 㥉���m�9Vk��N�ǹa���}Pdԩ��ln�����aӯ����N��̾8��� ��t�	H��È\�\k>�&���yB�:��ɨ#�}k�z�ǭ\<��w�F}7D�)�0J��Cp��#5'�m�&Q�Sne ��|pP����0Q�#�Wq��Y�֘����v�.@���uYf	��7y�!2^�F��\�XP���i�FhG��݊�YU�����ȭQ�o�)���0��it���o���^7��>�,Y�I�]�����l��+ƺ�^Z��T��;�(�[E�E�E��tEbW�O�;��s��"}���ĸ�Op��~�f�q�X=7It]�:=-`�� �F*�]#�nVǋ��$	`jq9�Ւ�n�c����"9�x���:"��a]�V��HGQЍA��KM5S���Ң�J?�>�;�ۓE˩Hf��v���-3��=rH�f�A��������&U/�o%t�[�&b�O�w�Ȟ����m}��)�sx@��+���:��%���R�AN����"����V`��x�ũ��5QƄwt�L�w�#7����;�5D	���a��S�oՔ��غ$W9b�?�����	�C1X�+M8��8���7k�� �H%��۱��ط�Ϸ�Ռ4
5�3դU`��H�y���wz@�wy�-_�"9,�qg�6�,�c��Y�e�7����r�ߝ~�޾U{d��V��7� 2v�J��ps�� ���_S ex}��4�����Ϫ� �'��ZT�c�#�ݎ�P��6���?��$�؀[��5���E�Lz��3� mv�X���N���r������Փz1V}x�ϗ5�����O�X���I���lJ���g�K���D��m�/�t���²�fr�ŮF�/|}��ȳ�	MB�vU���'�߄���7DZ/��}�B|�2���ŭY�.o>�������'`Z��e�oF�?�VX�k���y�?�4y:K�����q@��ߨ.�}1�v�d��Sn���g����y&I�����e'>���Q�X�R\f�\��pc9w���70��ނ��\G��������y1�Z*�Xv���f#��gv����M�,�Vz�f���8���&�9�4rr������9�vP����Ι������դ�Ql?Y>|��������0L釤I8N=nO;v�<��ư �"SR�8)EY�P1|`Y�ڬ���N����'�aQ���
lI�V��d�E|z"�P��DR����\{]���{C�����	j���;�yt�5�h�v]S���N����{��6����T�fA�v����"�����&|k�9�#[�`8���A?E�$M���<^}]HV�r�i�d�:�����F�K��q��_�_3�9~-��̩��}8�ԺL#�kW��=���[k�_����S���=k�Fc�d6���L��D8 �-��TI%b+�o�?If��#�R���ud��U,6�P���P}fƃ���-@4�GV�S��=�OjHTa��.��&�K��~äp�خ��-����tF�6$V�g!��ݨ�.��H��i���{����m.��j3<��h�/1'쯍�"v���x���7��4�D��^����-2���5�N5�h("-���(�y��%��z3֒r�豩�.�Y}�M� �j>})���qU/\�'<��cx�5�!�4���i�R;V�dTz6��!s�]�������ϼ�p��MפlA��H�����([Y�5M��h��&��9�W�ߦ8�v��%�U��+57�A�p�����pi��t�����ĺ_�t��=�R��@���tAE�r096.]�@+�>ԕ���}���q?iJ^���a�i�[>��LR#����OE9K�쪶��gfå_D0F���,A���[v����2�vZE�C� �9��E���1nC�d�M�+��p5���}I��c	UJy�H�[q���?DMѻ&�^%z�kH�N�=/|�A�W�S:�W���ؗ^T���-)�쪑j	����|w���������/hr*^�dev$&��~U���\$���'�w7�jT���_y����0a�+���3#�Ԁ�?$N�7h'�˲��T� Ҥ~�k�fVl�+!�hm���F����{*�*�����K�S�ڌ����K ���W\�>M��z��!��Q�葝)YO�\�Ϲ��@�@��w����Ǫ��O��J�%��$�5��ׄ�����-�4����[�з��R4Y�&�MDҙS�X���^Fݔ!DN���/�_M_�:�8>?0��K��*bvKLHD�t�F���-���E�?2�{�i�������������S�:��-~�em��Pd�޴�e����nbI~�ͣ��I<�|&��O����_��(�_o�933�����=�bL�ݹ�O�$��s��mnv��2 ���`��O��^�0Lm��_�y���q�Y=e>}ܝ���O���^�&�m�+!�h�Ͽ��o�Gby3�U4Q8�FHU�aq�|ʧ��?=ޜ�?�Ej����ܒur��c~��W-�l��w��PQ��'n[SJ��!���5.�S~j��o=���{�ɷH���y<������ǣd�m,Ϸ�]�����M�����߽0-�(�v�v�%�=mʹ�ȏ��Z[�<h�z?檕M�ѣ��ߴS.̷��1ſ	 k�<���-�����K��~�w���_��{���fkv�B�>V�cd	$�U��}A?�~���>~��B7��|۲���~O��Q?ʢ��hB�V1��2;L�F"��?>�ݛl�����J��\��5���Գ��,��id%=)�X���j��}�s���	� �J�3�W
���%K���e��Ok�O��{'�:�*6��,�f�jP��js�Qo��Z���b��[��(<�t}���s��o����Ío�tzM5��KL����~�����|/��{��7���`o�$1<oc��V<k��K���]���a�JV��G�m�&���@
~q����%F8��ޓ�O�g޲�p�穈]����	�u�=�QĀ#��}�Ҽ�B�#3����u�SX��ep>�d�8�g���]G��.ć?��sj��a}�c��G=i��5jK�a�]9���%:�R5�����r��ؿ��R2�q����Z���ꁓ��9�5�j�}�i��'���+{TA�o�9��!��������᧙$�j����o�f�D֢�nE#����o��/��Ņ�B���3/ǘ����:��C�V���C_W{��K���t���9�u佨\�;J�;��k8823�(ϙ~,��6�n(���U�q,=�3:�C�0�4�I��г7�ƂP^�K���\/\�	p���'�.����PQ�����HQ�ʰhQ�<�q'��xCܵ��݉-u���M���}2�ݼ?L	�M��Q�-3�7sL��G��n��1�JνN�.�{m�!o.�d�3EE5=����r�)x��^�=���;9�7���cuܾͧ7r�_W+X�=Si������|޻!��<nOT�����#%��I9!�ܶ��\���2x�q�K]����r������{t{��.��-����,��ɹ������|��?'�C�[����c�T��D�!w^u�PH��V������Q�\��sי-;�C��� ��),��EG�n�W��گK�ː�;)n}��o^_K7����{5p���7�u��QnN���.�wlv���l�fR�Q�z.��6���/���� �����0;'w%97ћ�q.DĚ��L춾 *�Zvһ�`c����勡|i[�tC�ڄ��陙�E���f��5��Q>֣�'Jj���NT�^����=�iJ��6���V|�Ac��6���g�qҵ���N�Ǔ���$���4%fmY浌��m	��G�gI.�NCE���<7G�$�v�?�\�^��==2B/y���G�>��i�a.#�7ս�
e�yt���?�1���p��k�)��o��g�)���1����{�Nc;NP%�h锷?�d.nb4S�e�����L���-\��M�`s�G���Ӌ����š���ny��ٛ�_qLi�ſ��b�Z>�� ̂�l�|�E�>Ϣ��D���BO��S^>6����I׃���o�<�U.�F�,`B�j����o�u9�����y-���噇<���4��a!����n������k��.��BFeS}�K�~����SC,.Jk���?�s�z�'�ְक़��e�
��SG+�K/FW�d��V�*Ķ��Z�{��䔽�uG��s7��W��D���L*G'7Az�Jn��Z�б���^֮y��=���`^�b�y���i_���E6~�̔=�����m�	�J΍�i݄��9��Y� ��ǎ̯�bN#�P}�:���ot�2m|׻VC���(����=��vn��t��&ԗ���V�7-`����7�������W@E�>�()� Hw�* �H��tw�����t��H��"ݹ�ҹKw�.����{\Ϟ=.wfޙ�yf��{3藄����l�I>���k[i��f;#�H����� �M�
G��!��h�?��j�*](�ۻ����_.�Z��沊4�:��&@����I�f)(�r �����҂U֌�\�]��;��k� �$�l��|�O˖(�^|z��Il$K����1_?�.eXȆI��+RH�Ҙж~�7)�t�6F�`�:�����Q͇���en[ba?�ʡ��>�GW_�����d��/�H�[׋	zN�Ҥ�OC��P�&��'M��\6���B�Bkc�;Kq�,����<�Ϻ���`�w�%�ц�h��Nٟ-1�7��ۍ�cͻ�v~ 9�P��8�i'ñ����̟U��\�"�OJ�r�br�m��ߖG�E�6� ��J��7�.�s��*�"VJ��5����hRf��z�k�������T#�C��s��&�^���?(#/c���1���+��6��!ls���-���]��i��������ܚ��#�;uV��k2��Դ����u(�
�[˵����ǶX��muD���S��rT�5�w�ѩ��L�0�;�y�ʟ\�6d�X���-��"wm�G�1/�g�gZp�d�*a1����t�k�m�K����ɹ����5ҿx%�F�z������y�l�a�8�A�M˿	�#�9Ҋ׿g�E+��ϊ���(슰�.�7�_�.9��������䮳i��?j�Q)��+�����6iu&OP`�F6A��Ɣ[F���O=jϛ�3�;�oz6�?��Ǉ����ga�
�nP���0�y#�sC���ʅ��Ͽ3��|�%�O^��H�K�$���"�d��?��Ѷ1(ߤ	E��|>�����q�卟-}랖���?���D�V1e�˻��d���٘�-eQ��7�)�QT�p�|��節��,�$�:��
�e��盧Y;{y#ǐ]�Q��̼a�]�`cVxZ���X�������Q�f���B������c��Nm��؅����`Q���i.T�iԄ��RD���}���Aر� ����I�tr7��R#y��g4\~�i���D��`H�l�2�Js�T�#c5�W�Oٴ�� .X*��Ao^�M��P���Q�f~ �N��z�� S�v���6��0.��~u*o�Y�?�H���ʪF���=tJ_����_L���v�'4	�-���^]�É�
z�RH�=�;�����e�#�?�l��C�U����n��6�e��	7�'�԰�3���{"m�u���c�j^>Ѵ�=������j�kY�7
�qn{C
�7F�歶ܶ���{l��CyU�@?A跆�
*ie�-���#07�^e���N���<JT!ɘ��`Jȫ"���	��aB2)�!��Q_�qS�_��a����F���ב!bA���qWʷF,��=w��jv����[*�a��g�':���ה�����W,`#�ِz�����A���J��u��dw� ���ꚟ��|?RQ��iop%�X��P'��L�k7STA�S�͵��m�uaWY��ʥ�")u2�ה# �O"3漈��Ǖm( �=��w'�(�A���쐌��D:�?���D�Ġ�� �eEo��Q�x�.�4e�0�DK$$�c�d�5c��f8���(MS��l9��l>H��s9WjB^��A���DA��*i!�v�o��[#V�et��_�:���{հ�~u�#�xy��j+�����󧊐�����q����r.�1kP\8���m�T]\,HM\�ȷ�brE�+&W��3?&��G��Q��7&���˗O't]k��1����,o�*5��P�?��c*��/���WZJ/rlTu����%�r��E�o����Hh����1��?[��j����)��+�� �K��aO<�j�����;���Oi7M�A���h���|��a.�MTh��PjL�q�D|n���%�u�Z�>�����6�v��>2������ířJYt^�x,�(��kF� �S�@6�F��X{	Ɯ�4��3�	��{���8� X�S����2�!X�򊆳����G`*��ZqzO*�v�"��:\}�g ց����ö�p��Q��0�+eU�(B_�N�&4�XU�y���	E�!~0m�v��U��Eq���"�oó�=��W%�a�w���*T�;(Q�1�d邭wG�B/�7������.w9�G��|e�Wk2�*�UƷs�h��y�BA׭7�C{��aI�yQ��e��[ŗ�3�7?�ݟ��npS�8K�nVD����GT�薉W�C���[?��I/9w����Xj��76�PVR�YA*�;H������Mp���9iЮv��z�Q��5/ؙ�Z���L� ���Pk��#� �� [%��d6K�?�]��v�l��7���t� ��߷g���
ǁEѸ´�}1�����(��)5a|�;���8N[q��u�0��S�0R|/{��i�ԃBWH��OҦ:�q��Z1t�i{(�
�զs��~�5=��1�lG�!��-eu�+sb�A@#�k��iL�V��P�Wa������J�k�}�e���6Y'��T\�	&4�������ņ:��agջ�|��� ���v�l���?UU�Hؔ|!�])���l:���M�yIϩ�F�������
!K��{�" �
)E�"�+�I3 �+&f�S.�
�m+��n����CQzC�dc��ݟ�w�f�m���8��,�v�	cӐ^/�NZ�sL(�����~��!�N[��H�llC��ݟ��A*���S�^����3��ʜ���
1k�����~˛H�ˮ��J l�e��l?���x wX)���\��}n�+��x܄/-M��k�o�����U���AB�V���LG5�9άՕ\ <�*����XX+%a�Y��ks��ek�\��G6 :M��!�d��1֗����i{CV9�'p롕}��"�w_�-9K&�]!vj��o3�`��|�yA��ђ�_ '��kL��l�ai�k�����M���x�� ��؜jVc�������I�մ�!�Y��̏X�W_��#��T���W�8#�g��~�-T���;�L��-�[�P{��#]�`#�N��(��S75���a�3��j{�ʝ�V(�lE#Iw�M��RQ��b���5�r��9��ǃ���grM?AR5���R�4߾��=P:Z��f/������~�zM�N�4��N�Z��'��a�>VY�K�7���vUCM���Y�t0A����}�3XPy
���Jy�l;�xAo��w��U�ɓC^�/�q/��3��X��r��ߞ5C�gy
���)��h3�å3UP��׭��!��6G)"6�]�2'�:��j�Fk@��ބ�0�p����#�ڒ�19��V6������Kp��U@v�4o���tP��Y����nlZ�>"��`y�3`[��������Y�0���ͺ�U��6��*=ɉV%�X�3���ݏ�S�ӶLJ�69�Bx��;�����_P�F-�VT��#\�z��W�b��@*x~�`��v'?\�oVc���2��Ό`m���j��t@��>=�Y�p�E�f5W��*3+E`�`8������*�����D�[pt�~P��d����!�Q#�98xQ`�K�>ʼ�����ߒ��݃^Rj�]��^o�����S<=�Czogy&�&��Lp���4nX,3���࠾"T�HѰ��"6���C��o��2�~�Ӄ\;�!r��ԿȌY~�z�BEW��]]E�׾/�]J8�)ֲ�X��sǉk���;�"�.�$�层��1Ȋ��|��d�Sʾ��2�&�V��{E�#_�^�{�B_�S�4����R��i�v�+�4�u�|>%ew��vI�d�~�e
�`���q�!;�g�횼۠����I�/L�+�����|[�*Nnl��O��G��FFVg����fZ��a�������amk�,����0��aJ�bN�� ︾��m��d�I]=��9����}�і<���Q�V������:"��n[SQ���O�7<�E�	kYgbp� Y�v�h���o�@<�+����>���Q5��]_��x�������fW�n�N��~�Wv��¹^6&Yz����~�U�@a��v�igr���~=c�\ o�S�-2갛0i}�6�}���^9��ix?mÒ��F��;ҷ�V/��P�;GA����)
k�ڮ /���?Lc�����ŧWs��z{�����(a�1�t!�Xҧ�����[�H����&�|���F���	�e�<uȳ.�U?��a
|٫�"ET��5l�v�e{���yuѵJ��¾S�vUv��d�%`])9?���`�_��Ī�<�_��Q6a(��Z����kv��Z���Ú� 8Y=w��6+��I�Q[K����.pQ�9j2>wþ4.}�J=��w#K�r3V{� �j�wJ%����JH�AA	�M��P��K��c�+�ZK��c��?+���.[,�n�2.�䩿����a��^���O���4�f�5=ŵ,s��
�~��ߤ�/�'BO	*N�����j�E:�S����P�����31�Y�������C����B�n�Ϊ�������jMӇSA�o��c�$	_���*�:�O_�7"moRl//���=][BW������D���(|��1YՂ��~i�/���|�%��8��91-L��=ۻ�Т���c7��gƬ������1�S�e�r�/P��רo���Uf�����(t�ޭh�C׳�$#�Ѱ�s�Ym���vR����1���Į�#�{����4���&O��V$~� ��Q�躤���[������*U�Mh��b���Ě;�Ov��!?��E��D�$��q�n�7����K���6�@�$Ӂ[A����^����Rjo�7�3;�a$i\�?J���o#ѻY`���';B!��C���� �D� &r�i�mky�M��/qOL�P�B��Q�8j�����X�7��/$rA��;�sƙ��}4_�^HL�"������n�)O>5�9'�?2�=lE�^����e�.��#(�5�����
������d�=ˀ�xnu�	T!foRS\�2�E ���U��op2����%4��O�B�lu���u�QY��]�yyh4� ��y��Vn��!$)�+R��Hа!��J3�������/7�n��P���#���I��U����'3np�e���ee��_3�$�0�YYU9��JCwR�y��⼑�q�l��Aj�h�ġ��k�R�q=͐��( -X�z��$���\/�MT�|�>�����郦s����1h���'�P&����f���ͩ��G�MDH&����'5ݱI���ׂ?_�B��C>�&���܍�%�1v�(l~x��7ғ����ک���{�u���W�l��KH�8��ʈ�e#�ÚL$ݿ-���~z8vp㷝vEY������.��ɕ|2���w< �4��ð���XH���pZZ�8m-I�ņ��_�KK���OU�8��[/�IEɋ�(
4�z~p�3��˼��B<! /�9rN��83^SE����'p��C{��4�����Fn Ȍ6�~�w���s���%Ue����(���U�?+n�~�y7�D�U*B�` �΍f�-R�"(������+����[{m�q&'�w��ZE���'3|U��6H�����9�|RT#��dP�ɖT��6ݧ� y�lGt*S*���4��2�DH}�sחH�
����������Q�j ����d��ggeu2��C�7��Su��>�7��EF*��%/9�.�V�q�NJX1l>>�U�� |E�V���g�Ƌ�/�;�қ0#���ݜƝT�νG۩C"L���8�dv:���R��
����߭X����M�"�Z�Y�>VV	i�]��g�G8�Y��gGF-zu��(�2��x�I����q��.m<����	�b����V��|f��&,��07:������G���0 ̯��OI!�C�6�2��}o������OI~��(�./v&��t���p��9�ý�ܬ�H9;I�Vp��Ċ@UN����(R�L����� Zr=���Rr��^���ǌr�1�h������7�5�;3��3+�d��R��,�7��W��燫��s9 )nW�Vr����^W��`u�
��B�֔/��0��7b3��*�,@t�|���nv}/���ۙ�% �Ʈ
ɓ�&7ަ�㈌E��3�FEW��d������X��*ŏ��}< v]B��L�����m�i>�l[���.�(�#���`$�~�����>��gf��$U�� ^� ��0�z\���)�1�P�<%�'-a����o&Vi�-дI���S5Q��ɛ[�}���GSM41��֟�-h�%X�MD��.IkW�Z�U�ɦ��2>�4.��8M������I1�D �[�H/�fCMJ��O"�<F��+7F��b�0ܺ�G0'��$�$�9*ȉ�U�rہ�d�xe��)�JI{ח�h�,6����L;��d�2= �������;Ԝ�&z�V����m�$���e�Cu8{�Rϻ<�+7'��Lš�8�����nc���������g��b��^Qd�4���V��B����$�@���k��ldȢ���7Կ:�ԦS�pv����r��jh�_O���������aWr��!Es"T��/[S�?Y��(��QF����h�{������:Hm��y%"�_+f믻�}����L>%�3�)�=�Bϲ�=�1v%1���ۑ�i�/wo�#��;�U_yh�|�y�_h�����S� ���J���bp��(ҹ̣�U*������Y�ն��1|������g�G1����/fuHv<�H����(3HI|���ژ�m�����t�cZ��2(c�[��7��cy���R��o	�&��Ƽ!��B���.f��~��
+(ޠ�%N6�@K�z6�y���6m+��"�C�A8�{���%��𳎛b-R�K ��ѻ��*���j�H5�\�4�K`y�X��3<g��!7UD�_n��w���~�vwY��G�	��?�q�ʏ~<�6dŋ��:K+�1����F�Z��ܯ��
��2,z&;'�r�\�EX�4�U�Φ=t�~ػs�n�R�����jI��/�
ԪE��]�~�)��‖�G?LW^z[~��Vu�z�
#v3��d���Z�U[���M��MWa<e3L�p�c��du��&��
����߳����*R�[�4�&�ƨ�����ch���ά�<����M�M. l&��7^�ͤ�ռ�f��CYQ�m�ҷ���%��?�4��~�w�@a�"ax0A� ��XL#����1��:�Tb��WC��g���@�y����I��d]Q!7��S�����jW&cV��?�NJ�ny})���ēP�D���5��M��Wg������ٳO��C�n���m7�B@X|'���}3�QZ�@H��],>�3֖�͝���*�&���������h���d� ��ï���"�G����Ы��v�fw7z���`DZ�WÈ��%:��Ȳ_��c����DQ.����rD���"/���'�0sl2����������ag�ДW��,&�d4���g��Pc�w�K��=�xy:�8̓uZ�&���[*�
����-�H�����՞wGa��'�"ހt�������=��#N�nY��æv�ew�羛Ԉ3An�&;j��G����IC�,��4��"�ע��^�k�@��Kܗ�k��Sl��B��e6�H"~O��2㇖b@l^���c�9+F.��~�MoI��AH��~J��t~<�q���ny�s���m[�X Dl�������]�OCb�Cv��{��{���M&����U�k�2=����k�_�N�cv�ǣr�y�g�Vp�҇,��ry�B��0\�>�[9�~�P���4F7��ɿ�|���M]Z��r�[� ��;�7Ïi�6��ae�=�3�)�ݦ�Ϫ%VK0��XEhK�o���+�2a��=���{ըĲ�z(Rf�Aƒ"HXm�^�w,�L�jA�qg�q}W��O"_��5�~,�@�-I7�i�ԁ��B�I%M�g�\A�k�x��aD�Eȳ��|�~��8I��e}�n�t�hb?k�[��u
���\�-��A$=�eۗf5��=;�Ƌ8�y"Gmj�#$�S�tP{�����]l�<�������Y��':��A��1�O�~^�6c�uu������$`tl �axx��m�Y8�ħ�R�I�vg�Y�k;����P1k��:˴%�"ѳ�?K�������6�~@�R�*0���M������j-ֳ�BV���^|>�V���5|T,�OQ�Q;�t��Z���0��ę]�y;7>e��E�]��C�4tG�
'��I7����Si��Z{��l��\:�o�+�C�v��]��5)����nG&Mo^��;��&'"��_ \��Q�O�Vv"��l��8zx�=�����;cLn�ko�~�!a��A���8��7�@}�g4�\�3�,b�J;��4F��<�<S��{]-!a�>pi=|��|Դ�9F�l�5d=U���!T��������~�N,�m�땦���#  ��
�EB�v(���k���P	Y���Z���ɥ�ȉ��3O�d����������+z�D����s���f=��׮_�}��T�zx3Q1��PV����5S� ���Qh��忭P��O���Y�	�b�eR���v�m��9�w�o/��Zz4孩�'��/��hdB�Q^����D'k�h�m\^`�N�4$ o�����u�\�*L�	����Lq����*��8�M�O�E��ۺ�Q����"��qP�W��Y���3��� �A�Kh��m���G�u�ϵR�GĚ�KU��a��!��W�>��'��K���=�i!%�� ����ъ5g-�`�g���sh��1��D~\�r�-ֽfu^����9�W�L(l5ȯDz�é�I/c�E�JFG̕�> ��hK�vK���m�oۢ��\�59h�^Α�1y���IM̿1���96֫ifv{L���Z�
��\��df��g����v�O&�k��'M���ݶХ@)����S	�8�����Lz�G`͢� ?&���� �* �;NB���b��6�J�+�p��n'+�]�q��)��Y�zL������ U����q�a�5$ !�� Q��GX�u�Nq��|O^�Nn)��T�^�����sX�M��{r�rLW�Ӎ�{F�Q�5j�<�����Ƨ���*��]}�<����j�I]�Ѣ��"Wۺ� @�d=~\��8������yz7��'pjt�FV�\�7<�e���-Qw�F�}��_T=̺ۀ�ҙ�ؓ�]{���?��<O,���Ħ�q��0�k���u�:�d��$ۭ=M1� l.�����d�.\���¡��r-��1�~R����$PȻ�z��(JK���ITx���=���(V�OeX��i�_3�⎛�Y�N��MTZ�-P3xr�R�Gvi*|��M	L[lMva�
&{9х�����rv�mp�U��=k�뻐�=E#����e�,K���ϩ���0n���mQ0�����j�М�:�6�����Κ�!a΍ǚ����P���?2���+x��O��+�d��h|X��f~��J���[��9^����Ӵ,��MdL�� B�0pP�PhԀ�S�d?�廡V�`k�i]��`����0��8�<̎钨>x.�@�@�	�нR[�Y���^/�G"�����;N*K�E��Q�&��( �BwR�h�Ģq�5�M3+ �T/�/�1�|� ��wY7�/���'�|�)O��0d�57�$�|��6��� �Nv1/Q��z{6(�bU�a�t�t��Թ���?7+��V�S:�| z�L���������c��4�5�<bۦS�'�d�͘.X�C�dzQ���]�~��+�,�4#U�WnB���&2�<^�'�\�I��_TJ�Dڈ��el�dϦ������$����$PL0�l��	~�T��/���q)p�ϝTl���積�ڳk���	�p�K��ߑ���{���N�N��)+ǟ<M{�<�jDÓ)��k��aO,��X��nE�O6'�t�X���ң#�/���R�F��8]�)�J��['���X)<
��kv�*�z�II7��w�QhNL�h���>@�J�r���y���ſT���+�n�>G��
���=5��h�c�9���1Pr�m�~.�R�-J#I��!+|{�ߌ�6�:�i�ن�p��5��קW\a>�E�'���Q��eŜ�ڋ����K�Q6�\UJ����v����-d}8I���4����c鬕��S�n�Lc�T#�f+nqt�t0Wn�q߼�i$}Cr�'����m8Rh��c
�
�@"!7Xu*h	�D��{yi�J�N���{�v���&�3��K�V����<0�Y�Lr�F�a�Cq�f$M�ӏ���,��ZV�TU*Ƣ[\.�՚�c��ȧT�*f���\��z��1k��d��
�Jj*_��ԛ�
d�d?<�zTP��̎��ke��K]��U�PhN$Tf�m��(|�Z]���XuYQ5�^/�I�jێ��;�l����G���E풌8��XBJ�����"kEj`q�Lp�ߩ�p���bA~bOk}�%���T�3,�o�Ig���g���g�E�����59\����(�9��x_!��^��[h�j��R)<���e�� ߔ~���p뗏�����߮�4��a�:gDh��t��c�����o!�̷���Yܭ�F.��ʙ�W����o�%6q�?���B���u}-�-���a�vz���2K�
5���S�7l�f}df�ݭ�@#ә[�+l4��X��:�1�:<���0��c�7�8��:�]{���I��/^"���Wn����N�r�'JRïg2��Č�L�N[:����$�,7��-�up��Oo���ش�WN��l
7--�^��26|q��L�V�Jq�X<��5S�x�,����Ƞo��3*f�Ә'����ɭjNX�u#!��Sߣi.X���L��+X�ׅ5��t}�к�nV߫�@թ^3���a���B4���'���D��e���ԇ�b�Z��e7�卹5�� ��25&ǂd�P�u��c�?��>�)ɕ�J��`����Q\>�g�{��4��M���o�/&���,o���	i�����K��a�
��_�4[����ܡ�Y��D��,u�m���v�b�K��+`�tb�8���=f=���H5L����0.�0�Ӥ>��	x��/{�Z��L-��n;?���}�p5R��K4��5��b�D��|Zr�t���d�? {!,y<ĉ]OǣKF׭3�xU�HMg)�u��5�ߌ�ף<�e�W�l��cr���
W��@�V7��1y8�,���y��-�����lb��{H��ߌ��Ū=�ȫ1�Zk�$@[��rȊӦ¢��7�t�P��Z�
��r�@΍A�(|���;��C0�&��z��쨻�U�.��$��W�[?�E���z�� ��?�i�K�3�P�'n�_��� ��y���H��6�>�G�)��l�N��0��lX�Pu�d�-Ȓ����A^|��ۺ-E�� ~���Z����L�0�'�X���і1�H�̤�X˶�w��Fک� ��Y�ib4a�7���-���
��g8Z}~)ѝf��e36ב��'���5� ��D���Q�㌍d�V8`����T�Z[�����O2���輪���FM�M�����"�������_g��w��dN�u��P���5{��;׬�Nlvc��@	?���I���.IҶ��%�ra�S��_�v�R�u?�k����ZD��р6��4�y��/W��B2*<��#UsH�5�����fЧ�Y��LIWp��"H'xv�>_�$�n���,l�&������m��v���j3Z80���f�r�ޤ��B_
,6J
������C�����#d�j������ᓕv�	9M �exY0��͜]ޛ����fm�j�IJ�%c@�ӆ>�j�i�7+�^���sx�^�-�G��(�Nk�k��J����x�maT[2)�/w��[��C/vD���^���T�:|4��x��`7�J ����Ym�jAV����C�Ut�T˭e�47���/���[j�-���]W�I,2T��K��L��B�=w9U�d��������L���Bq-�Zב����;��aSq�/>���J?�p��I��4����B#�Iy�'�;{D&@.�'���I:�����c�r�����mְj���6�ǲ�![n�(T�$�
͢OMS�	+R&��䱶�~���^��[����}-���fV���f/�0�뾥�IQdV��|r!ޜ�x~��gO��q9��+Bg­�\Iu�,'�Gw@
ɸ��J�8m���Y����G��'���}he�C��L�C]�.�+�6�
5��`aOv��N���w�7��i6�5���"�sen2�@8&��+�c�L���WueҸ�����7�e��֎�w`L�ơ�\Ԁ�t1W��}�l�"�v�m�:K�y^��2�y��6I_�J�~`��e�lqO9����|]kƁ���Y��.3f�X�m\J��"�0��,`�#�t�ӝ��^�	��5�B�����j�$T�w�����~F�&|	y_�6nm���.� gRszI�� 
��kf�j�>J����­
Qe�Wxh���o��Э��H�Yn�Ꚛ��|_�:?����t�}���|R�d1%�~{1&yZn�G� ��fm�@�͟��<3�U �{��(���h�,�J��1���f��b���\���.��'�����	���cx쌉��a�B���`>��F��`��@��SV1���rq�h
:����Juj���ܯ�т⎔_��y��@o'�@j�p���S�}�w�� �s�Nj؈sn�cƔ�
�v�g��|5F>b����h�,ZY�5Vl��k��|���|���,-�ļi�w;�q�Qf�#���k>�맏��g�2�R�"�g�) ��ّN�w7�����|���#I�$8^�t7���� x������w�N�t��y^�Ӷx����X����۠f�FH�j+��Mr����ß���C�kQ�T`=�?wO���
���}L9Oe�泸0_0��lu��%�������PI�1�n]��s-[ �i��9\jj��^�1�wr{����dPk�!+D���y�zr���+�O|!��&Lq�s�i>�w$Ԛ\z�GY�J�b��G�V6�P�$"{8�Z�P�j5�8:��f�j-K��\�J5�Y�oh 6�m<�s�-�4�r�gϫlg�mО�ScF���M��P��:_�I���L|�)g��7�hw�fsm�u�����s��) �d���S�a�ޥ\����;��J�����I��x����zS�%Ł��I#��)���y>��N���
�N-і}��?�q`"������L�m��f}��1�� Cr�H��}1����������oI�	�W��W�_��~���K��o�j��P֪�pW������F��\�f�_�B]�ܬ�w�Z�T��w��V�=I�^-I,��T��x#�{�q���,�ۻ���K!���_r�׈��$�'7�@�:������0L�	��j_��������"7�sd�Y�h�9�)�� *L�(�(�ON�GO�o��2D��C��;�}ҋ˭�������`֟7!z֕;�T��$Ǚk��f ��!�� W;�߇�u^{j׻�;�d`:^��$�����;<��q���%��c����3�{
�᪣w�bS3&��y�B��;o��^\��եܠ`�6YB��n�_ݖ�ר�8�C<���<�.���)*���咏E�R�A\��T5�L��S	K︕�]:����n���Yg��_�7�٨�!kH���E���L��v�Gd��)i, ��5��1p�֙�Z�%1We�xJP(�NjJ��{nN�Z��ǥ>8��:bg���`&�I!N��Vؤ���pD�[xf|��p��Օo��i�~�����G[L��U|�3���^�`�f�-Ӓ@���N��<�/-t����X�Fs}�/�::�b�n�}�Խ�>�85��tG�c�4�����|٤[j�s� ��۬U᡾,���������1MoNg��'R��/��j�A��ϙ����e���� �ٓ� �O��ɓ�FԷ6{�A�"G���|�g��;Տ�:]؅��/�2$L]#j���<��_OV��.��{����4Go�"�l�$]°Ļh�t@t�����"x	b�w>-���?�i��j,�c"�L�-���`�}\G������a\m��D={��>v���w�H�cTi\�61���{}�.�VR���2M���u/W��l�wl�芛��>:��6zBީQ��l`&-o�e��:����>Cf�*^���2)�\[b�ˉrg�y�0�&��_n�8�5#{���ݶ6>]D"��&۬?�Ť"���ϩ��n'_���{J�#����D<�D$CKnv�s^7(�Ĭ�z���D�t�eD�4n8sc�u�h\����T��(����4��p��cc����S�o	�87�>��ѿ3�*8��4H�=�
�#��p��(��A��.S��y�$d[P1m~�?;�h��B=/�$�Գ)��PH����dr���M&�ՒT�`IB���?�Ȓ;��g���裞6�(o�M����yK�T����Ek|Z��E��w�II�JL�����%T!�I�}ضLS��6gGs���<s��t�L�x杏��n<�?`[s�5Fo��y������-e!Gy)qk����p�L���iJp�"��h��F���ߪ�Z���k��&�T1�٣���t���0�~赜��ǩ����г�
��{�i9
�-��ܳq}�H5���^Ѿ�E��?����o�k��T/�m��Y�^�M~�����Ǘt4�V���;p������ ��ٿ)�*�aZ�w��`1��f+�,�s��0����X���c���C"i=�6��y��b��f��r��J��{S��o��6j�ㆹ@lR$s��tҿE���M�X�$�gr��o�j���n<ˬ�!�F�}t�K��uJD�5������JO���݊��8�kSϚ���/�u�ql[�84�N�f\�]����z=�y�i6:�/�N	r�)P�*��W�	Վ)��u�ΕrJM�Z��3D9�d��5 Xn��ț�$?���u�(���G���AOك��(�lQ�_�]����z�ޜ!P�oS�g�K�����E��ֶY)o�Z� �Ԙ�'VnbĮW� �M�d�Jؠ�ʾ:FʢȆ�2tggPRiG�k$U59dna�8A�+�7�W�9��|PYe��!(MoJ��z7�-K<�O�A��鸡w" ��)��"���:��Y'|y=�H�I`ȏ�O� ���C��T���!�<
�o�7��)'��/�]�����ܞ��O��(����G��F�
bܽ3h��{	�t����Y� �0C�������{�D@6&G���_NaA��2�:��"�;�/�A^�\��[� ��s�p�_5����؍U���k�.���dg�	��d�Y}N�/�<�m|߆�4�*j��jW�o�K��p����<�����2ߤ��Z����ٛ��4��x.\�k�t��]b�}"IbՌ�M�r���b���Mg�>���\�a�3^�D�/��<��\Es:lNjaK�"�w��hp�A��1*�x��ۥ�ã�ַ��}N�h����5�Mxqξ�;�R9��e�e��d4,���B205D>؜�M�a�ӹ����Uv��5���4pC_��=���;��q�6�=[g̜$\W���� �����
	����u�6+K���H2�l	�23�B]�����|�L#gy�Ʒ�X
��b�er+3�É���H����j�&�(�)�KH�q ��[@�怙ܾt�l=%�lc�c���X_)6�����X�tgD	;�-����kMk� :���BDO����@y�@�	��_�&O���~�7�S�����xC5����¨|�o���
l*�o��w�o�����6mh�_!/3Bq�w_�q�\m�bf�[�l�\�È��=�w�뤌�&�l� �����pw�iՏ
/º��v[} �Ů�8�Q��X8�@8$�h=qw����.Zf7��1��$_�%��$9�N	��j$B�Z6��^�������� Z�l��8�˄깯c���NP���J��_O1Q����k�Ч�L�CW��?Kgr��&Ó��A�l��	����h�u��ɩ�u0 N�\;�~��J����5k�w��EP�� -?T�~�8&��X����w#�6�h��۫���L5�f'%�����7�2BJ����}~�%E��)��_n~�j��Z�$	��Q|����Gq�&���̃����:��zIXO����*��ή���&=��Bf;���37І3���P֛_ :6�;ᬇI��5v�|Z���ЭM ���^��G�4ۙ�M,���}�<ϴQW�C��H� =z�7���ؿ��r�y���F�F�^�z���J)p�%	�ME^��{�ay�������Eq�'du�D�ڙ����j���!�釲�F�� 4}����wni~n�l�٭�%�oO�Q/:Suyb�:���_ǘ���	0�>��wY,tYU��0�GQd�0�g�����
�&����J�EABT�$%�A����Α�AE@I���k���" Lr��n��������\�5�s�s�s?�s?��<ȣ�);@ůӯ4I�R����k��=��{����J�H5�՗(�<M�q�w8e=��^��~h3d��Q4��'Ȏ�/��0���~��{a����l��� �����I����������q�~qj�((�B�N���)eP՘s/���l�6��)ы�3�nt��T���T����t7��A9kgz�9�ګǟN�v����GsxE���kmЙ�!h�s�q�PsC�ܡM�D��feF؉��l}�5�X,��5+��x׃I��Z�Y�J>qbKv�C����T���K�X3���ː�3�1��'�Z�[�;�{en�ݫ����9~�5E�ij��M�t!.D
��i�tJ�|v�j�ż@�!��Z5G�1�,ļ�� ���{K/Y�����y9�ߚ��ܧ~k�Na��u�
����IA�O���tjLR}jV-4e���}�$%��t�^sXSq��4(������)���bq뒑��~�S6s�M�K��u#\�*�-����I�ⴱh5���P�d���܄�|���A+������R�ue�#����:l�r���J�UO|P����t;^��/n���x�c0���Z5q�ո]6��gI4d������9A��1n�߸�?Nţߩi��� l^0���+�A\aB�LCp�5���M�uE�7]�?�Q?|��g�ib��K�ި��h���^e�*ذ:�R��dC4�ks����
��sWy'�����k*O����3ˋ{b�V�9?��k��y��R��ˊ"_F������e��F������ȢY��Q�W[h_����ox���KTZ�-� �ma��[��ߜ����iT��:9m����I(���D)�y��p�'�1�	c����][�|�S��}����ϟ�F��<�T޳��4��G\�;� �4+�3��TСP���tU�|R2����������iF�&�4k8�_rͰ}�T��n��0l����O�Mo8��҄Y����%�^��aX��a���W��BE;���.��a�ְ4�[��ȆF�XX�m���K��e�8����������Y�\/v�(m�kd��#�~%�']P���m_��GtS=�:�qP��x�
譟հ�(i��m�1W�}�Ѭg@Ȫ�{pO!�=�L8��,�N� �2I�#W�ܚ�I	��`C��� O|!y����G�i��t�XHL��.f	A>}����{"Zw$��O�j�����;�D||���؏�!s�L7�,C�L�6�P�
���_�������gse3�@`?�i�>q{ǹ�S���L�h�Q
��� �km�QM�V��AsZ�)ҍx6_��x�/�Ș�G��Z �!h;�2�q~6����~CQ�O��$�16�?�[?�F��@߰�N�@q�|ȴ�a���@���F�*U�FU[��%݄ "j��*Qp���mΣru��
�l����Y��}�旾��
~����N�8Z| ��X���GN\�����L�!��=1�n}�y��A�X��CIS�"vcJ[���T]�R:����O$��U�7[EeX�s�( 6�ӅH����g0���"L�g�����ѳ��pjn|���8S���}��N�\F�V�,~~"v65*�^غ�u,��>tKo4[�RA�eB�C�N��JJ�?�0��(E�D�E�s��6�\��|M:!8�v��g�H7�τf��PD���L���y'hF{nm�<�b��7���M�F*�CO-dP;F�h4��'�R�¶Kv�1��������
��^/�K{��~dkb�6�0���X2�����P��<�O�@�`��U ��8��J5�,Vy6�������X�mܔ}GT��D��5i������@VlQH�H�n&�������)�?��c?�V=m��}�ɾ8��A�Y��I<�io������Q���|��8ä��{?�:u�0h��_%V�)����?:��ج׭�>��9l�BG_����V��]�p�C,m<6�r
�sz���i����`�O[�����c��/���H=88�f}O���

歚���;��	bn�QD�5��%�l��_N�����`�C��l�ƒ��e��?S�6wGr�	�hF�����k�C6A�x�h<�xv6~8ee��d����2져����w���+���鎖��ke^Oye�BQh���M�J���ky/�K�͍kS斉%G�ڊ�N�dp��F�����m?� �}f�[`{��Q�Q��2���!|O���hRc/v���ܹXS�&�'���~��^�[Ŝ����~&gg0�n\���Ay؅	 ��H���'cD��^������>Q�
�?e��M�Vg�4��]� X���xTj��9Y��`JDө��l��q�<R��'y��G�	%R��T�?.���]ށ'~oB7���_X��'�ŝ��~�	�p�����L����=N���0q��TUUGY�^�
}hr��Y��Jb�s-5btlynܵ.�YW��%E���&�:�������`85/9�`!�g�;�^]�2�!k4Y��-��PN`��e�rk�s�L+}Ҭ���]sJEwaV�����l `��G������������q.��4�3�Q?���>�6��l��di��\Ɲ�Df��F{��:�b��yu��܂N)o�a�g�m������7��5o�����jy{�� v{[ޣ?�~�z���ǘ2�e�?������PZj���N6!�S�H������[�N��V�|�'�8u����_D=���7�r<��M���儎EX�_��� ����ω<m�m3ˎ���L� ����d��N��'�d�`c�=1��L7 <=��(U$����h��_��jB�C.Z�Zu*��<�pT4Q�:�hB	eS�0E���E�#afIA$5;	Al�hS=����A�@_���X9�<ĄY�[�h�(B��Ukܻ~}e��B?�VNJN�9A��
+�mLtN��Ʀ8�xƧb��a>��S����2SPWu��U&i�4!�_YE��#�J�J������g�aN��]��^�le	�!�1.����][������P�k�C��L�@��������rӘUy&����<Ys���P��B�XZB|��7mxa-����:�#��o���O�@�������`ޖv��C�E̰>��΢�=����'oO:�,iu>0!H�-ּ��\xDo�'��`�:���Y�`7����Vs�Rޒm�G���D�+����摄������s��򓤺��a��Z�qN��{�R���l��nR?��0S�j�k��tz�gT�J��BH�'���oǧ����4{��U&�70E�ƫYv��Tf��a�h��~w���'Ɠ��T9T{��&OM��3�bi�[=�w���Y�.�\����� �u�ynZ7Ρ���1Er��&3B�/ڿk9�%e�G�!M�'7����#��<Ծ3za���ة�� !�ka���ʓ��##�i���{���-�����4���L�㔛����;��cv߹Slэ&r � �o@�B7J����vyG���S���k��7w<W8�<������/<�cai�|&����9�ɝ@�N� �p�]�)������zݽ�E����)����8Ό�h��v�R���Z0�p�v�;�V3�,��y�R��1���[�߿����p�j���Cb\�C�΋mt�!q���
��N�Z�^����녒� 0a�U�G&��?�'@Na��}Ί��^�uܤo����_ܸ1;Y鋓�fX�����s>n�����X�Fc��m�7�t�R���R�4�rw5��C��ř�Kz�^�!�Ĺ݄�H��G�]5b�%[��1��g�?�pl,>)&6�ߢWC4�Kؿ3��+�EnG�{��N}�����o���k�����8Ojt^i۬	?\�H�|�-̍@M���u^���k�j;��j��P�q�h�A0���|S*m��p;��uC�$��3gS ��e�Y+-Q`��C%&=�X��x�
4�+n�`�ώ7������&BE���T����&� ���'��#e$Wz���0�V��J�FI�(�Ѳ��/��Z��D�u���_^��;<�e-��*_he)�^�YE��S��^U�����ʈR�&��vxӣ�Ns<Ȯ��+���n���JT���y6���k��<N݆�=fK_���N�#���Us���r7��@#���ɥԝJ�_�N���~	xQ`�
���ˍ�oY�R��Qp�q��~v���Mf���Ѧr�>Bd�zCt�Y��Bݦg�~�0��~��R]6�E��,uX�M�b���aG�jΉ�p㗼��o���[�u~�%:�
�Y�%4~���sLt��C��Fݣ�fC M�<����ӣpǶ@ў&W�?��^ۚ�rJ������}�61t��4��{�&��XKvm�����
����F�%5�[m�~�M6���AN/�Ƴ�8\��&u���^o�\��;c���5���D
۞���k�8����f��3�=VK/|F��EX7T	����U;��|1�b>޸�i��yk{@��6�(>7q^@�.S.8�������!���~���I��^tn<���{�p����w	$���e��2�Z��D��!I���3^�F�2��3��@:C����u#��˞[��C�0��$�_UA1�i�_ZbD�AUǧs���KM3�������j�}]�ܖ���=�憩{E���?���7�����_i?��Q��ӉM����{V�q@���C�mo/���/'�D��˸ ��$Z�?����'/�3�"�`��e��J����=^����?3|jD~A&�����<�d	�y�ƻkO_n^�)���g�e�=N
!`%���k� �a�醲{QY���� �� �����ѩ�,��W!�cm������#Q�NJ��Y���O7�l��m����l������c�gk7O|l��n�ے(���~M`����A�������W��G	��]~#I�r\B�ˬ�NH�qω��5�Կ)8N�T�[C	��+����H_���M�W��Uf�Ӯ�^ؚ��\lE<m���'dGܹ��v��w�w��<� '�#���bƗ��ѠNx}ه��R�=K��jD[tnz�o�Mt!l��%m(KC�b�JH��Jl�҆6/N�EF�&�����Dݞ�[�u��s�1rV�x���̿y�sݥc��� 30�Lm*�{��2�h]]��.�$�)uS>k��y��١�(��`K'���H���}�?���z�[?�m�o������ZT�<��8Ȕ�a%�5"I���O'�c=_:��U�|A��:B۰ǂo��JV��U��ޅ8'-W��|��+�m.���Vege2Uo��X��*�v	������7�|�v19NMSX�}�ST/Y.����9��<�hIY�^W ����.���t�S"S)�b��jq&l�#b3��woHl��z�	%e����{պ�lD �K�����?�`�i���&Kg�8�Ha��*r�%7��F~��N
�m(�����Mǆ���߽2駟;���[�o`�-��hM��ש�a�Afv/[Ak`/$_I����ۅ�o�s�w,���Sl��@��?[�;�8�@l���8D��z ބ�i�q#����F�w6�[ҺF�Y�,�Q�������:&�;Uc���|�@�7��R�{o{���@�G�O�wV/y*1���[N���3[�L8�sc;��D=s�z�+1���]�;��9�2�,D #R���G=+�.C����B��~B�GY0=P,lbj�[(�oeB��6�yؾ�4mrЁ���5S�]JJ�����MV�V�a��A�b���,����1!��j��m��$�%�����s>^.�V��KJmv�&����N/>��4���Mt���Ȟ�|�K��������ty1�4��Z��GA����֗�wq�O�|w��x޽'w^�x�w����s5�t�����m˛p�5ѣ*����~*��2G��<̧�������hKy���|��<�Y�K�X��dS�a�z�X�N1��Zyp�ԒЀ���
�9�k�����&�ּ�?���3�����ŕ�z��M��H��C�o��➮Ϊ3SP�㴊��_��J�W�f���DQs����F���1Ð��;�Oɺn��#�U~g絭�=m�y.�W���袤c&_v`SFS1�d��gjw�D�H2�"��i�AbFh
(�sn�t�9r�FQ�x"/�1�
⨽/s�5����<
Y� �ذ����R��8����'��5e�qX���d�����T@~[�pi{���)���Y0MoJ�,�9��bB���v���8Z�=#,��A��H �n��6Z�BM]�<�r"�K�z�>�"��ӹ�^g,ؑ�7�6~BBI3<���G{=��ۛ��X������/@����X�RjF�6�r�����C���V���R�g;q�օ1����aR�dԇR'u���G�D��p5���|�V=�O��lސM�U谐���f�0� 43мU��We�^]9��m�����L/�Wﾑ�w��&`�����6���I�Zw�������D󖰒��D1[�~y�N�Z�N�w�g�IVi�O��D����J+�/��,7_��x�2��}�o꺥�|�_H(�1_58)�*3Ū^H'��6�?�+�Ϡy�8�ã���:�jn���v����V���3��}X��ՈT�$2�0��?,�����iw����
��pBN٩Q��=bi��X�6�ґ�'w�EFa�3�ub�V�JJ�������_S�Q8���x��4�*V{ �����`�F����i9�y�����2
����'g��U���T�&6?"�;->G���Cr%��)C����TPj&j�*[%�b�\��[�|y�#IC8�LK�Aރì��j�Mo�&�8�� K΂W�HYc�ü�J�M�8�ݓO�"p�n���r�v~A�'�/����tK����["`�G�	�6Rr�-h�:|@r���!��R˸�G!����g��@��h���mB��ĒҤ2(�H'�dl�R20F�^OCi����u�c�5E�a�&=�<�Kwft.�"�z��>�9L�Y@-�(1���G�����HPXص�v �*�O0�tӛh(��n�R����H�E������e,�DjG�5���ɧ�*d�#�i�_%�5$�o�2����I(�����A˦GkMOL_6�
%���K�7M+?A�<բ{⊟)!"5qIC���p���ZuR�^�<ԄrϦ��n��L�~��%��d��(������&%G�P�_�:�~���aؠ;��kI%#zx0�ˣ�����2����\��1�F*z�^C�n��X�DTU��td���*P��Q#�_�9�(ri�����l�z¤�]W�#���4Y>B��x�T�����s�W��b���y���EV$�}`�Xz��-M'xE8W!�3�5䮔��y�T�=�y����x�	b;jݥh��AtOJ�bƻt�'z�|�A)X9=�� }�3N-�"B2�/�u��J5��`���q��(�v�4��"����枱6w@>�0��@�X}���E�W�ϭ����*�R��t�X���N�\�;�
�Iz�=[�L׺��X���U�:Hbjۜ�l�"�l�?"���o/@g��Ss�3��*d�,症�Eۂ�D��sg��U ƚ4ȡ/+:�,μ�ݦ� -bT�O}N�u�xU\�X�M�d�M�GU-�j��w�_:�|��"�>��L��$V�31l=����,�fb�ߡ�*����� ��M�}��x������~�{b�f�c�~�����f����҂X��Q]o��
)��	��Y{��3�M�jY4|]QwO�{��R���8�̲tV�����zh�;��v�1��]��V܊��0�����?��-׉����#>]�_l<z�"�0}���h'�9�n��ϐ�#1	ɞ+��<��V4N⽍a���UQ�tG�(���H�הZ�6��+���yy(s�@�J����SgޫN\�.��*<�T 5�|&h���G�cJ��-��k[O>"�jݏ��z�y�kS��U����!;��O;1�!�o,��.�wY�Qu1Op���Pֿ|y|��ݘ��^���j��s��g(Q�z�2�������;a�LH�E��=[�5�x�4y	uJ0OT}�b�p���gM3�6�vU�.��q^�w1;pnKײ����V�Q�:����& lރo \Z���C��������p���ZuP�8�D�7�
o`�]PE��ٝf�s�n���v�+N�!6�)�Ey�6�9ž�[�Tu(e﬎�Q0/�-r��2�����]}fn�!�5��� ˟/�x/�������?k��"yH�^���uZ*P6�����Q-Opm��xZ��A^rF��U'��� ڮ3zK��/ͬȝk]*�g�D3
���\��Vtھ��Ɲ$�"5D�Z_DH��I���HH�~.mr;��ߛ�V��P�����3�n��j��$KN\��}{ f^ 
Ǯ>y����p#U1���0� ��t��L��N�*��_���מ2���뵻�S��v]��QC�"�\G9̞���V���,����k7 \�8��H��A��Tj�<��xL��X�έK�y%�t�)?/Ya�d'y�xX�B�ާ �CѴ�+�T��R�2����T�����"���p�eA/Y<#t�����!ٴJ���d�r7�_��k�
�P ���]*XlS����3b38)���p�B�J�5ĢR�a�+�;,�n�X'=����7<���z��PGI��9��_l�Z�p�z�XL	TTn2���uQ}���Z$\�Uw�C��a��PXwT���q�V;��͛��	bQ¹�$q�VHpV��~�K�c�喅;�wὪ�x+#�y������w��z�r�qC�I��n�~��ۺF�Aޢ}��g�q,�F�nIy��\�� �_�|�sn4�R���S��Nq1�ub��1ǽ�s+�W&y�Ǭ#��ɣ�v�'��-)Q,R�L�����Ǧ�_xfv�� a�Y9�������۾'�R���`�/�%��b{�"�#�v��m(�^��$�6fa�������x�-0��F��G��/�c�ʪJ9�1�P�8��$>(��[v�B�Zi��c}^��z�X�Z~X�J���J䍞�=���<ݞ8�:����g����y�ɜS�bõ���%ou��*�p���r�jy�#�XQ�{1�գ��J�������nCz+�de��қR��lx}�a�X9�yu��9J�m�i�d��}��y�1�g� ��b�e.�` �l�y��S/��pPy�g�h�n��՗�skL����R��GZ��	�9J���N<����}������f������N�"�D�6���/h}��
��
)ٴxZ�W�w_Y�:�ĚdE�.���~^$�|ʰ�������ݞ_Փ��.8�gѳ�Yi/�E�W��`��E2lS�a�$�[�w�[-{�����6Jm��ᇳa#�
����ڳ����Kߠ�X�R��l����e�ɣ9d!g�����a��cǐ��"CL{&����e� b&�@�*�������B���q���ɾ��P�.𚊑v��РQ�+�$��T�Ğ��O�����.OܨD��M���s����|)������@ō�@֡�b(=�*=���8�\�Vq=�0l5�s�9�}��K͎T�
ѵ�§уD�:I*�K�.�jJ5sЅ��'%�|�a�,u�{mM��C�����[8Z��2KZ]7@�@`����v��;j��\aq+�IEO8�^��K]��Smឈ���O�&s�vru�e�������sEd�使��	?�R^]=���c/�O�fř��`�*EA:\V_���^�6��5)&o����Y�*ϋ4�[S����fI�L�_��8���$چ��m���d�:-	;y9�L��J�Q�OR���y$ߞ���U��~W{lpT�f}�\tyB��k(�z\��S ���w&^˷N�ک�-oz��$J?+��ۇN��H�%K�:I��1�W/��4���NOg܅U[�o����E���t���.v+�>�6�����*����V�P8�$��և33�itH:<���8Ή��YB- ��i��.rr��R�+��WkE��r�VZ?�c+�	^s���p�͜g�hk2��AڟnvuM�C5^7���.$�4_�B��k��$���`b����*-n���?W�Oݥ�wr�{��u�w��;�m\ҝɜq	��z�w.ʹܘ_�;L�>��`����{�&���aK�B�ӛmeK����I]e��Ip��aE��n��˚���\�]T���]��������S�@s�B�#�R�{���oh�Se�2uۀ'U�+1����s�rf	����A�8K�|(�"��ñ:��c�'6i�� �Y�c$1�<�IѾ���A˄�uR���w���]���l��1�[�9R')t���$h[D~��+W���W��0ʰ\�@6�cVw���6��a��x�zi���<�.�ˆ",��.��V�,�H��� ��9��!j�ލ�?_\�#�7e�b�i��Q��$�R��U��2HS!{+�
�L��[I��{8�@�\�?���_�x�����O6<����Ry�kY����9�S��ÛϜ
�ֶ�ȫ����N��ep���S�������eG�v�!Sj�a��=���Q��D]~(����ҽ�}��-T(��E�9�ѰdSP����X�7�ҏar_ku�k0��O߲�&-�.�)s|r�kp��,9��A�=���ӥ����rK�[ޠ*N�l���|�Pm���C����})
�YG��c��]T	OHS��6ڜ�n���d�ޞ��3%T'_�i�|��2���1�.�mF��d"K��h"�����L���yM�R
k�+8���s��sf��HI�Y�|�t������֜"4
sƺZIz�MR��߱N�����~�H�[^:�;?����>u#r�2�Cs�����4�DÄkuir7��!m£���ѹ�:�L�K�{b��0�Ș�߶��*�ؗ|ھ�&�-���S���W�I�Ê��'�v�w|S�"�MD&�����c�*�>O� ���%b���2�
Y��V��Ƅ}�4����yֵ(����.�����ko��g<D$
�z�SV�h[��x;�<�"V>�ȧk
�p�W�N}ڀcT��&l������7_m�ª����.o���d��B]���\o�*ſ+E��a*���D��P�ž@1�F�(&M!5́rk�_��ћ�	�0{�1.�L,�?�R)�[��^�% ���)Nx��Y�p��p�\���x�*t�ħx|�Kǯ�?"�~EG�ljO����j=*���;X�|�_3J$J��佔�	�Z�,��h%���+��Y�]��.Z��uA�I��˂���6Ź�k��8@%ZG��M�C�C�70*m�ح�`�b��ש�k@�L+���Z��A0s?X�?F%'�b�/yM��'���3Ƽ�Pgp|�c�-�f��b������X��N=mw|�BVծU�GH�1>����GY��!�?��%�������������H�hHn\iY\D���<�_X^�[?���l}��b<�?�ͿBՑօkl�`+k˻���٥��-�!4p����,.\+}kغ�����ϸ�)�z�Q�+�2��送�{~�?�I�D�mn�wV��If����݆8r�+��7c�B�B�dp %(Ͷ*�3��`Г>.�A$=�Kx�إb�Я�aG]V.�cSwVU��X����4�qFT& +��'9� ��/�.t��%B�����;�|�V�3Y\f|�y����'M��7M��(�}���Ol�e��effa�~��}Q>_�������l齃U㭯E/��a�#����������۩0˞�յ��r%�\jO�� K�l�J����M�Â���I�hvD�PHVoZ�� �
#�qym�%�3����A뗬�3�u--�R �8���,�ߚ���A7,b�pa��As�O4�C�	f������(\��k���-�2�?g-�:s�JHIy�c#�=��XL�ed��q��p�K��q�<�vՆ��O�W�����L�U(Ye�9A��
�]����e`�\c�Lfk��&��/�7C�b���Ў���ݯ*�~�w��ե��Nr.�sYcqZZ
wc#aU�7�����S�ږ��{#|��,̊���䕉Dĉ���K��O�n)��/}*��IL��+�c�ǔ�~<�3���>e�-�ǈ�z�|?	�y��*���н}u�)H�4�(�z򈂁�����{�'
߁������e�����a֏g��������Z� �;��vĨ���*�^T��������!�?�Ζ:)����>��������<���h�<�I���$� �|�t��̪���>Y�~��]��u�ŃiZ��H���������>��,�N��F�=�G*l��1t4�����5���nW-#q��~uYlv��9���J����|N���Ҝ�['�d�퍶v��g��Z9��΍��s�FHV��B�T.t��ΐm˔.�4SJ;�r��g�K{v���]�ۥ�}�I����U�mS�W��ߞ���9d�ث��a<����>zy'K�g2�X����]����q�U�}B���2	S!�)�#ϵ�A��v�8i5K�%�m}zu�	�s֢�q���qI�Ԍ��B�?�i���'�;�t�~[�OLstYzUfK��V�a|�B���In�؈��A4�����[�?�<��,}��d�s�H-�)��'�!�@	���럚\LF6�F9�=�h9���5��V���$(���J��k�2X�����v�6Kxt�D4�<��n}�O怳����&Y��>W�T�L[Ssdb"��ނ%%���.���~�X�����v�ڈ"���#�IEcr����9<��i�v'��D�%�ջ��y��b�ㅏ�>*`*{��Ϊ�t��5�,v�+dWe��^��U4��G��.]����J�A��0�;C͕���������L���Z�';�W6��Y{�o��U�[u�k�$:L��O�})n@v��?�=*�;ݗbYY㦸!-�Ӕ����!����*���7�̑��p�X�*�6��T�u�7{�}�9���Zǯ���������[��݅P؈��B	.�D�ΐ������9���d4
�N� ��G�v�c�����`�+K|g�@!�>��*[R�0M�zDI�7|�K��t��RJ��$z�K������~c���K��A�ܩf&���K�Sa����u�'�3ś��K�W�|����d�AY۱�RJ���(uC+ nA��������\g��k����/y����OgP|W6{���_�M�ۈ)w�x��&8)�L2�DX;��#j��O6���Z��/� ��2N8��*?��\����$�PJ�k��̢$��a��+��)	�k�U�����q+rv����驏��Z��uk�i0��u��pRT1G5�xI7�*��Q�_�'S]�#ʿ+^|L%���l]�����e�?y�C��ӽ���5Uꪴ+���K3|��#J����=!�����H.eb�k`6/`�M5&m"`pF�����,G�ɕ�Wk��3B9��sɖV���1�>w~�jVD5�) g�Ř����B��!�q	������l�o ��^������M�Ð�4nE/DoZ9�Ĵt~��ۥI�-J���k~�����N�{���ى_�[�ro��G_����b�{�������L�j(A�4�nr\�.�=࢓�ž{��.d�_�tkbFΤ�B���N�Ї��,+��M���+J�5���x��AƊU�B���w�o�9�>C�Ml�>M�(��|��+<:�ùP�7��ٸ��YBe�+D�?������sʾf��M�!�Vc�z�#m�B�h *ע��ɳ���?��ϖ�Ò¥[:��a;��a5ҖCL_�S�~�_�=�#�Ǐ-XN�W���Q��.\�;�����m��]�����oKw=v��N�=�e�MU���z2����ݺ����\����Ý���d�fL���d675��Լ���fV���DL��2�\/�:�%�=i�����=1��4�3F-�j�7�L�L�`:w��}�L~y����ɺ�nr����t[�_� -�l�	�u~���sgi��h�#���5#h�ٲ�u�H��=H�:�o��j���djW�S�^�Қt*yQ��#O�|
�x��ED>|G�A�&����T�I����W0hu�q����7Ơs�9�*�`}b�IM��4���T��-~��|di*��E}��=�\����&�n[�ʛ�\$�oH��Em��f����C=��#Ak!R���Op83�
��x�d=��4��F0�ǻ:�*q��B���o]՝.��%��e_�٭8�����<gw6��>#<8a�>1-/��Y�
�g�
hl��<D�hE:+ �]�Z,<�64z'��"�#A���ݝ��h�c�cH/F��R���<�.�j@h5o�]��*E�I'���.L��?g �16߽�f�����P�\�:�cZ�;�®˒�?=���;�
Rï<ʁ���ϸ��������@����Ē���mb}&������Og���V��ua��	ZL������G��3������xu�e��c��j��6ҁ�!�o�UF���5�Cb������wm�Nܮ�D[KHܡ���
����	�p]�@�2F	�m%�	k�~]�H/�_莗wm�45h�H�ni�f䢊����sQ�3$��\��G6`<�ˁD�����dm�.�����m���2�k��&��6��A��L�.��r�@	M�B�b �<��}R�.���N�;�A�&�_�����V/�L����dI��PU/0��o/��1�7��Nc�m��.�U!	j�=U��H�`'y��r	B�Gh}�ڪ�K\�!j�� $IuC����j���I����dߓJ7t���6	���Z}
�u�5fb�F<㪸�]��k�����XG��w�#F�깚�
M���N����ͨ��A��Ir�6��H�0j�S�;E���!�y�g��:��YY�O��E{es�0�6�j�����̝��[�O����I/n kU��M-w�#ϼ�J�� .+n��?Ҭ����Sy��:
���}�Ժ9���$���?Sx*���~���q%��,W+8$��i��?v�Z�v�k9�Xs�4���}�(�=`����R&�1QN�;��GZ�4x�iA��8�%����O�7��`1�0��t������V5��7�4�P@��l?Ǒ��@�_F��L�+t�t��.�Y��ΛzD�B����i�?�7�ÊJ3܊��K�h���vF�̙&0��d1; �(PV��O�~�kW��Ax_Ѽ��E�����Ȑ���=V
^����+_flO����r�^3�q���Q��]V��n|Vk*m�񲻨BoD����M�ݯ��Ռe��hhh��TEz���N�;�<&�-��Ҟ�����3m�)�
S���D���Y����I.B ۗ���62��4�~�*t��^�i�?�'k�z[y�b�:Ǔ�~F�竡�ݜ~�6Ƽ�pŭ�{NuDn�&gJ���,���|�`ei]xx�a�u��Jd�#�K���G>�و�QRY[�헜�����@���~_z�5��?+l��&��J� 9�1u�	p	B�J��PY����?�S��"�p㭢��l���%��S�AR�;�fw��O6�)W5��ui�O�(�Kp�*����W�׽a�j_}�D|����qv�1	�to*;�1���x��}�ҪY酯�D�D��'����	fUy^�OcD�P\���;��Q@b%�5\���W�:��dR,p�GZ� �x��)�yUr�]7���+���#q���x�[Щ����B2�m�*Hg�֪�l�I�����t��o���cX�Ũ�}.�y<���im{pc�vգ��7�)�:kU�Qث7ɣ����|%;�ؗqK��Omq�
����jZ��#���f��(�8�l}��	��v�2�H�\�=\���ϔ�K=��Ej��W��>��@�*c��"�H��4�XrPJkn���<��-P�N1{ª����N�ۏy�q������Zi���2qtI��}3*rdc��/IɿK����m+o�V����/
����=�%�b��y&��vu�H���Ck�/�	��8���y�e��$H�`!�LK�����W_����NO|�ʴDV�q�&To�!Y��������C&��JN��-��".��Lh���YQ��%��o�!����x�8�V���<4�d�#9Z1+�������Ur�=w�s1�z�un����WG��n�NL�f���;��f�;(I��K9���U�z%m��8���
z5EMc��p�t.sd~�R->1�sGJxOIpo�qn�?2�~���N��/���l�i��l��@}+� y�^BmM�h�z�������H�6�����F�f\�kM1)l�$��G��O\�(�SǶG�K��<�]Y��(��6@br��$�B�����$��.h��ߌC��z4�Ŷn�������1�i���o�m��̪�����5ްo���'�����!"|��8���5`��r��!g�dېdc� ��T����ո(��ϻ�t4���q�Z`�Ы��o�dy�Cא_��L���x�c	���~�T�uX���>�r��4��E@Zb@Z>8t7���I)i���Ai�������~�0p��{]�1��콟��u�{���d�����L���7�����PY�o���S)�;�`Q9�09x&��Y����%�p�ay��Ur?��,͜�3��~Pu&Ǧm�=Q�\po1��5f�I�7��~���ޥ��+gqrݚ���{�%_@�6�n��̪�ܡ�V+AZ+o����X�$\��j����V,/�$��2 &Y���~�保Oy=�h���ߐ5��>�(� �q�Gq�M,,�a�i��{����kZ���H�0�Oee~��r���Im�Ɗ���bl���Y���bB���wU�6��T/�é<*+y�)�H͞����t����3�F�-�?����a�'�2�*��rS��6e���)Q�[��FH�5�~�]B����j�[�u,R����'�2��5�9����y$��ϝ�
]rq�˓SṂ�9 ��~�O�$�������Q�0 ��~�c����A���ΙYY�q#�>��-q�^���:��n��{?̴��6�����60����Sp�������D}I_�>�k8C?^]w���--Tu[t�(�5�˷C3�>��\��@lё�8�$]�縧Ɯ ����@�緩��Y�㒀�r��^�����f��,�w�"m��`ך�gC��C4s��� }��w�u�Ǥ�H��3�<8$"SX���ɑ�yΨ��L�/5CU&Rp�V�q��>�g/*;���}b����=C~��|$��������"��yͻ6�_�q�pok��a��|_��dW�9����>�j~dX�_]H�]����C�v?��z� /�M������ �,J��|����y��HJ���G=�,�`�r����`x�Ȣ�=��Q/v�D:-�����ыgv��/�Y�yg�Jw+����e�������eF�6�bO���m����"�k�]cGݏ|�oҗ���:~U��1�4Q2�6��<�z��>z� �\}{��>�?�/��8��9��{��1�Pp�9h�W�uQ�'���J�{��K5a8���&��Q"Zs��*MTs�Y��9Ւ9:�/�j�٫;���Z�0���	ͩ��@��ُ5�>Kd�3ZG��5���OW�����3Ym�g.�ۖ36`���2-ȏ�l���.j�t������MƓO�'%0���@��zf���Z!�"v��&�0���6�� V�v�mW����^κ�����h�	�������]+�_ӽj���mYAO���nw��M�rF��4�ء���6�Ú��.&[���'P�tnQ=K#�u�S$�Ǵ�a����w|2���N�Z��_�Ӏ@M���`����qn��
�����}y�;sή�F s�l����WSy� �%�m�
�ͼV��I�`x���k�7�[6٢����D=��c�h%.F08�_�H��u�J)/��R�I�'ڝ|�3��Y�\X%��_��d5lp�۸�|c.�z�\|�6u�x���TNjw�l�޾����v�M�	x�|3���dz��I�q쏧�&��Í�B7"��ji
R;�g�
KL%m�U�����a�ө�Ɩ�����)��2ߢ�a�1r�OA���[��65�g��I�zYuK��/`y�0,a��ZO�Eh�H�4��&��`��"�p����oj/&�Voy�1���|���k��;��+�#�Y��6�]?̈rF���㶵.g.�J�sij���[^�k*�0�ӐV=e/�N&W:2�d��(�~���qu��X�XprV$h/�%�s��!�\}nXU�5o����X"/x��`�x_���Ǆ&�_V���I� A֢֮2�ѫ��.�2Qm7��р\b�0"Y��D��N���{��5#��t��N�b�!ѿP�"���r&�H_��~ȧ|�GP9�,��O��o�&�?�Nkz4�U���oVZ��*)T���{�m�T�ٟ,Ud}o1�k_ ��E~��t%{��1�W����5.�����5ܓA���O�u�Ň�[5�Ø���-�Z�Dy����GA���s#�D���#!%���}Z`��[���STs���3�]AX�M]"�=�"�*y���A��	r�'!*���x����6ɬ����ٽ�~Aĸ#xr�d�u��5 ���i[�������!�t�E�%�!�n������������\,�-P���<_�
?[`3d�r�J��2bm$ 2\�r#�:���$ǂ�e9ʉ�+��@�m���Խ�ؑoG4>+�f�05��xˎ���o���{0\s��\��[U�x�*��i�b�D�Z4t�i	<��KLٶ't��zY%"4Qs�z���Q�k
_��n����]�����P;Ə���$���ik���-���2'S�-���!��kG�m+���9px
њ��%�(I�6���[���	.��k��sfzJ|U�a'�4i���Qa PV��	:�4�A�Ƭ�l
�y6��8��1���F�R"����e���Q�5�"RoR	-�g�ʤwdf|�I9`Z��eԳ=�@�Hc�Y��_�U����(m�5$�I��Z~����\}�y+�����Ȕ�o���,mL+$�0�a�R?�\��zhTِ��n�R��p��0�͙�M��$�S��.tJ��A���d�1S��O��;�}��s���軐��"B!m�
l����gR���Q���^g����ϔ�3=��sy�k�#�y �r�]��w/8�������	�2�l>l0fi�#4�~yN���7f9�QҨ���A��f��`e�	�ԛ��p�삢�\F�=� j�"ݟ�_��WG��>g�T���#M���|�^�Msᙒo�$.��c�������j���O�g-<^�j"��S���~�G��B𱯣G�א��N�G!����\;����>��7�ג�;ݸW,�%�>a�*���b͠�vfȼ����ݶ*��-V�/x���]�a�'h��f�M�d�6b�RA�3��az<�r3'��\7�7q1��ѽ�ԡ��.����5uٻ`�	���*yc�芚�2�)�%�G 
ٶ��5+�"��a�޺6���{�Ý�#�#DQ�98�E�%���%���C��*v�3�"��:"�T�j��eG���) 3}]�c�Z�M�������%���Xa���0�G'-Ӟ���8Ѩ��8:!�ν�eF��f�}%ߜ���QA������}A*�8*̂��;�*�h9�5� �
*�bv� �Ɣ������79���F#����Mw������g-Ж��]c���7' �x�l��D������j��'/�N�Zv�a�K���A�Ҙ���>$Ӽ�����w	�54�e���%�'�I�\y���)�Rq�ಣ&H?+>d�%�h����(�u���VV�8>9hF�f��DAEncv?�@g�]��I���غĤ�ʨjTfG4��hf�w(����wC$��CÂ=�5)dY;{�q�U�Wg>6��Y%zc�]���5)�BP�"@tߜzْ�yFig���Р��O.�d�"�h��ؒ �> �i�
LչMs�Y�(���|.�Uw�����ϵ@F\�w����-��$5�=.\4./C��ҳ���7�V�d'!�[�yV��2�H�L��"C3���Ȏ��j��9��&���I��#� �qAe�ַv:�6&vL�YH|æb)A�La�KX�^v�����i�6�)�ތ��5�o����]����^��AUlF4Ź�O���+wփ�h��?����h���C3��֞���d�j���˽����f��TKO''ƵQ�М�Ώ��ϙ�<EFC�`��|X�����2��}�]A���2�6�����ތ�Z�#�ӑA��~c|�O�"�x��pK7a��*��3Ws��N�.��@��4��4p򩋩����<q��k�����"�_tW�0��t>t˖�����FQ���·�6̙����M��d����~���:�K� �W+�tr���Y�����5U�|��N��
��`�����'�'W��:� H%ٛ�ڰ�τ�Q�������>7f4��'���_���$Ŷ�&5��a��@S�����s��`�\�+����A,��^��L�c�
F������T�S˛�:{8��׷�^��^�3`�`��B;��8iQ�Nt��x�P�<m����vaQvb�@�ug�:�|d�>&����Q�A�� }7�-�J8C�:��5�+�����yC�%��;A�X�e����͊L�I�ݐ@�#�J+�
1x�S˛��`�\�@q�J�p���Il*$��ypV���	����S�yv1�b��a��s���gi�+*���1��Ig�����u��@P�������o�J�/���[�t�p;oK��1�|'Ųa�������>��2�+S5�{DK=��J_��k*��mqfg�ֈ���X'N��&�d'��S2����/Yq�s=�3�S^�;-!ݓ7鬠of� �D�/�j���J�9rf�}O�:�T۔��	g�3�O���T7��V�b�.�1�$�-Zg|ܝ���CM�x�u�B�$VW}��3��oLF[hzR��UVk~�Ѹ�I^�ɜs,��B���8�8��������D�Yx�1����SK�G���T���k�T=4���s�ܣ.�#�aZs�̆B�,�{�*�E��&=:T'��#�Y�7j���U]����zO��XUH���C���'�����QSǲ�A�Ep!�ْ�J��W1�Suʍ���X�Ɣ\�ap��ze8�Pt2n$
��4!��X�Z��H��޸�>s�������U<�-����$NNS�+!�G������2����"���w�<zQg8t��{�;(�b�=WDf��U8d�ꐖ�kd�����؃������p�]M��J�V�E ������Ȳ�<���'>�zXT�.�����HCu�xw1��fd��$�l9]ubU߀ut��Y9��w��V��SXXM7���oD�DU-�Z���"�s��[��� �(.�Z	/�7r5U��k^�9��H���Y��c��a�������ND:}X�>�ցw >�+�����p��ⶅ���@�a1Ɩ� 6+��׌� ��5�i[��a���&Ph���t��zh߂��E��D���xz|�g�tTq�/��������s̚QR�P��ԅ}G�#��АA�T��p$i�p^>��WM7G�=l�.�-kN�lq�z;G7i-~�m��~k~>���!I=�ku�eg�	yb������|>��l������5��	��&�ɱ̱��oO���Aό38k��g�$9��n��P3v�����l��s�mQ����ګA�`���۩7� �N��̶x�:s�쐵~���ޜ0f��_b9�9�K� �
�a\��V��#��)� ۂO�R�\�A�1��T���i�{~,�v:;��#U�O�_������-�~}WQ.�&G����O�m��D�I-��I�Zsmv�-�����Ί���{��!.�yx�\
��i�[Eo/l�/]�.6���G��?�A�s}�ڥ5̽�]�T<t��h��7�0d�f�*ɰ4hµ�fҗ��ԡع��S�d-d
V��Uἂ���o�a=�RF#�P���L�<Kn�`�V���~��.eΓ��u��۲H$�~�)&7�x}��:/�>0J7��uaB� ���S��4 �|VFDjp`�D��e��0]e8*�������1�{d�����H�\��ͭ긁{~J�������lP�0e�,����D�Kd�"�-ʃ���:7g��X_7y<�1��3��SD[2��"�|�7$�o���܉0^��ڼ�s��={�L�@���7r�j�έ������U���9�����} i�Ah�&+l5���G��p�@wg�f�Il�Њ�ڢ��+E�9EoS�ݪT�K
ª?�MvQ7'�}��@y���Ug2��6^�A�8�����rP��k��饓g['�����"ֵ��Qg�r���]c6���a��.k�|�x��U�#>U�Ǜgoc�_79Q��}}�ˋ����yNr�!m�2��TNjց|W4��ޢcr��
� <"<[��.�Ng'��o��I'|*�����O$���|K\���NQ\jԥվ�#;Ra���[r���y���m#vK��d���9��']�_%<:�&m�s�>h$¯���>�.W�*+dEںy�r���*,�Ճ��hL]M
�GL�<Ts�<�_2�̊����Φ�cl��y��k�#g����V%'Dc�Q�^n{��$r�K#�`Ҽ�[�'V��	v�J���������.2?�G m�W�k���w:ZH�G����]�����(�+\��Yf�x��p>��X|�8]�ap�5? ���)Mv(�`:t�����nB�j���\�֒�[�w9�M��N�q�,j���eE��F!A Ryt��8�e���?��{L�Ԗ��=��Ƨ.g\6F]挓a�c�r	#�QT�pXP�.�QT��f��A���G>WMW��G&�&�kSr�"��J_L�����@�84��S��"�)b�0��y��{O�([ޡj.y����_��`��9s��S�D���I۔�Ծ�r.f��l_�xWA�g�R.
�۹��,�)@�@�U#<���N,��U9�zzl�"MnϥuQQ�Q�L����{�w�}�>�A��l*�rW�>��e/H�z_7�0�"aL�؟�<��������c`pe��b(j�����h�"��3̜u��V������٭�t(L"���e���p_NR���Y�y����� l�Cm����=_����m�0�]=�9�w4�d5`��z${�w��r�|����>��=M=E�WHQ��ɵ3���k�b���*�>�!h�E��s����CT�U�����A`�w3��L��X굜i���A:Yd'M*��"����dU��*/�j��}��Y�XLV0,�i/�����$[��݋��#���׾5v�L�w��~U����띢^���V� ���FV�:^��D4���P���mR&a�I���y��1�r���K�~�l��.<�25*���7��3�r��8����)�dq�XN�(Ԟk>R��M.ڳ�MM`c�o͂�F��	��u9�z����*�#jv{)C�]0n���"�����P���ݩl���EG�ݏ;U�i�3b,j�	v$���D�Pu��n1ŠK�2rn��ҵ��-�ˍ\�E0�B��p�B4�5���p��W^ѝ
t�7u#HT
۵L-U[^=K��Θ&HH^�B�z	H��y�|����I+�vj`+���=D�_���u�w&z���|g�0�}� t�|cl�kocӎX�����B�n����G8�D1�DD-���n���D�g?��6/&���E��np7�]�OK�~7���ɎH��&�uJ�i��,��GJ\,�MT�\��M�֋+��r��4N�m�Sv��'93���>�O��kqKZD��_��:"Sp倾D���Z�o�SOS��σURϣPU�P�zg����Յ}��$q��R?d8�;K\�#�?��	dF�`��Q��Q�i�������P^q��' �H���� �����z�:#�~��mw���v��EM�#5�{�[�d1%�b��?h7|�q� \`��R�d|�?�+7��۫5�G�����'��ݓ��O��>��]˻�����X��,=�Z���8��ˋ^�����).�Μ1p���l$v5�H�TQspY�����q��.�@g����QB|9S�m���"�����Z'��暟J+�1�-�Ը7jq���]�t*N���_]�:m(���J^��s��@;��q����#Zm����KZp�6h���s�4�~\>l�ށ��A	�ϻ��0X���IhB�����g�������w����0F�7:-ܝB�h��h�*�6ǉ�vW5ꔊ�/�F�d��I�C^�~�b9�G��%�E���p]�&��Eg����t��Cԛ��vʢNsNЩ&s3�峒� ��� �h�;F�sx\��Eƹ�	3�o�	�u>H��k8�	��{C�ms��9�rB6���M���/��G�W"��$6�V��~��kSѱ'K�o�:6Uc��dy���c�����VH������gI��N!�Y;W�=4+���r�Mp"܈��"���@?�=�����Fxt�?*����S��9 �t���U��n漓#j\�q���f��,�þ3�v��mx�'���P���rv��I��O�*H<"G	vY9b~~4�ymt�C��9�rz���a�Кm���5My�� ��_?�U5����1 �bd+�����D�LOq���� �Bv�4|kI���Z\S���j\��W�D��^����x�r����߱J�_��0.�A��f�إ�C��|�ڀ���W���V�Q�&}g��z�ј��m�-��Ҥ}��oj\�n^F���c��Z.o��[!q�l.�����()<R��[С��ۨ�keU~N��nT�8��αR�����?�na�O/7%�I��\u�PK����W���$��ޗ�_�dMX3Z�t۴I��񻄣���i[�|;����(8���q��a ���f��UKq�Ĕ_�eL{Š׮x��ob�Qq�n,������{�E	
���+�[���`}�+�^���e�#�����2��Ze�D/W!j��K�uA��1�q&����"��vt��Fx��Y�"tj	9�ף�I/����	qf|�|Ĺ]�����l4�ȫj����_A�'zT��`��w.~k����y6��d/�[rv=� ���Um�E0q�x���O�^�˟�_�m�/&� �%��ca>� �񨽲U��\s�ҥ�(�&}�i�0�yI�?]�A�"��q��b��ȳٞ�f�Ffۤ(H�K*N2��,���/N]$�oh%�.>�ݬXLS�J���
�-fZ]U�]�(�ڭ�����5="�X�xΪ�{��g?]nTg�J$\׾.��'��A#|��i��O�![Qշ�	ַPV����j��.B����>�k�:a�̳xC���wK������>�pĘ�%:�a\K�	MY��"���k�[G3dY�:;G&�韖U!`�\iv��O�""��6Y�n��h��1O��A�\.t����P[���P����6R�u]X���W�o�<�HȓJ�ʄ�,��)5����ڪ/M�GK��S�Ӈ�3����t�i\�nݕO�襉���x�i���S�J��K;Z�w���>�.TIܦd�>K�DK)������wG�<ђ@\W��L_hRt�3(��N��3L��z���s���$'�?
�m}�`����N��=�?h����� �����c4nK*���\F�J����^k{�c߼[����P� h1�_������}V�"����^��0�[r��n�%�g���)�o_c�v�{�ȇ����K���S�u^br�{.�ʷ�10����~�+���˭���8�;K�?��=�m��I�H��ß`>J�̼�Sy��>��JoVԶU�?(���B�Ol�� ��v�p5�@Q
:��Z.��,��zow�����XkE�T���	���\뎯�Di\�w*�|�v�=�.���Ĺ�J��~�A�Ït5l���3-�����8�����`�Xi�t
*K�y����).q���Ϊ������f�ɭ"4�'<�
�1���u1R,'Su��X�{ɋ��_�܄��R+r��5��=�ey���ݘ��Dh2zHuӏj�$t��`��[�?�%�K%�j�B]�;^�%��|�[��S�SD_Y��Tږ�+�~)�Qo�1��r�F;��2�9��i?��MO{)�=ޠ.p"�P�M�C|U1ss��íT4�+���6��O��"�)�z�jW�q]��Zi��4;��a��w?
N��V�$�.
�~���o�y&DJ珏n��Fx�M��gc�3��Go?�8����e���\�����Â����˸�����1�M<�l��D'?�4�F*\rT�W0��x��U�B2��6��{w� �����J�~�L7���WR��GL�(O��\��6.8�i*���x�#�]ß�#� ŵй2s�(ƞ��)�W��w�Hj�M��ӗYA�O��F
�φ]l+�>�ryZ\��je]��(�ku��O���*y��ٸ���g�ۮed*$�kR%r���U{�'T��*,�*P	y.���M�y_~%������Y�ɩ42/a��5�W"�����].����$�����E��ZL��^�8l��X戴�� �0o���,��� �T�TՁT��Ʀ�����;gM��I��Q�E�<�uH�]�!��R�ǤSZPf�yv��E�0sɺ�a"�دpt_{Ɩ�rm��6�KVh���u%}ݕEz(��Q
���/|=ƭݪ�B�+O[D-�n��>��6�N��k�o�z{z�Ϗ"�\�_&�L��Ų��g�2��F��}����B���V�2�j�ו'�ڌT�l�U���x����O���*h�r[-Y�l]�~���ɾ=+Q�&<�����i���X~�4� ��i�I'G�M"�m�g�
���0��?�ZZj���^����}|�R��Mc��j�����M�%i������nE+��w�F_$� =��[�\��E)����p�71d����u��?g���i=FY��{cW�[��oFdd�>�.�}/���(�����[y�mÃ��]�$��99Tޣd�+��w��/�7ͅ��<6QKfT^������I��#ȅ��GIl'��^�-�o����C�ru&vN�"CRٱQ��C�����QbM�-Ȳ�<�-^-��׾z��JӉ聢���cq~�~[jƴ=g�QA����D8�'���ٔ��5Q���5��N	)����8�1:L�P�]/xu������Z ���ѿ�_e�m�!<#C(`0��Y�����V#GYt{U�+�+�{\��ێX��(���u��*7~�.D���UX��-\0�]Û'~���k�e@ߛd�rf�/�5�a�"��Y��&xR6:1����&{��X.U��⩐�੏�b��7ow���"y��ʝ���ˮ�D�!�&����=g������d��������kcty>Y�Z�A����ȔT�_rA�%���{�2���B)epk_J��O��qɆ������oW6 �Iq|��t碗�3Hv'���{�z��D���������!�uY5�%�33��o��<8�v��kݵ����i�;̢@r�g[`����x=,S2���Z���nE4�V���:_��G�����BՆ�m/b�F�bJ�R<�כ�P/�υ�&�\#VE9���+�ZE8Ɠ�i]zw2�$9՗4���Xf-��$��~\�^R���4�&�N>47m���D����/6:�_̈"T(��XA:P\T�SeO����%�q���^�-����uo����or�`M��'J���#�%?6�~dS#�cW�}}��ަ��qF�H����!�Πּ`�
s�L�Ujy=�s��F�)�Aru@)��&34�����wOH
�k�AOA�Ӗ��n��4J��Gm4�Š�b��H�����QJ�0�S�*q�ޛ��������Oū�58}�|%����W��~�l�G~�VX��
UᣙOb���ǚ�):�!��y�p���"z�%�V�������Y7e�e�L��adGxB�O����u�M��� ���A֐�q�$����хA	��țj��x�J֣ʊզ94���!y�%��$�G��[�i�(J���i�3�u�]�.�t|DU���c^�Lë��DW��q5Bg�2�挢��j+V����ꋻ39��Rϸ��w��׌y�œ�'�en����Yd�PlV�v�3�5oi����,�MJ���;��0�.�}1��L�4ں��E2I)z<����_�G�Ob��@۷�.��IV�����nsJ��_��)��{�K~О�+j�Ľ������F�8t_aa,0�4���b�lñ^�l/�v�X\Į��Ԛ����Q��U5�x��7�{�59�_�{7�b��CFV�
�8��LX0�*�O��u:)5ꉠц�U��B"oݫ�z��Bo�$MX����zn��u���f]�'3�s��;}��H@���F������ڕ|�&Hp�$j����\:�����@b>{����eBטˤ62�2�
ʎ+�F,`�V���N���k��D�6 �gXY�U�O����ٚcO���H���>�i���g�t������u�l��#�*Ņ�e�B�����FS���%�A�;��u���@�ll��c�Z��3'���8BD!�Ǩȓ[ꃋD@��pW@� D�pwd7��>�`�wp+M����E���vj��>��Z�����30j=u�գM�a{<�ҟ�9R{����K���~�"<b/9ޯ�\%�%'(x���_P���t��b�"��l�0^��z�D�6�z��F��[�m�f7����zdN��J�:�5#���p��9ҥV� �*K�U@�ظ�HQ�1cO7�N��ƛ4�c�HA�l��ۏ����F�.N��ץ��i�?�ɋ���,�M���}�b�XU�D�y�{�7"2D��� ��ᮝ����@j-[5]{�ą��k�GM����Ή��'�6<��~m>$%�~�)IM���%�@
�#�.>1�.o�ˇH��)C�����u������S�+�R�k3!�Q7�4���?���v�M���� ͱ�W��Zi�Zy�#G$̹���_دӕ�7�0����w�<B*s�
r4 �ۼ\qq�/���,:|�oӍ\���)�,�~n-�ܟQ{�;G�Z�����y��&帉����Gq�W!�}{�|�zӛ7�d)i�w�9�~��1|��/��3g�)�!k���C�N�|'|�&��ͅ(3햄M�l�B:l��؄�xѠ�\��$A���<��%|P{�[��4��!Kc�wz�X��P�������Bi��nз�2]������o�~6'��nX��Wܝ��ř^>�X7��9��!�w��+�i����xi�7 -���6�1|>� Y���!F��݂��p�T���f!�*�2�j!��2 ��k�R���������ȧym�o^9���ۇ1��
��5��v��#9�o.�wE�i�-1t�eM�����DC��� �IMKS���Ǒ�/5�ب��"�q����M����:�F޺���E��F�f�v�*d�a:yZ �,���';;�>�2Qg2e�T}U�[BB���Y7$���צ���޴��u�� ҙ���ѵ��a�d#�MY��n�&V4]�z�j{�+,��pOr�R]d�9�3�
��WnX��؇�"�)�>�6�je���Z`1�@�*H�5��w������m��E"���u�,bj8�����`�P�p��Y��VQ��?7z��hs���p>�Ǧ~���y�E�vW����B�&lXY|���}���c�5�{P��OO� Cvrz5�������/#s5n��Z��Y�����F����-��0�]p�8���������
�U�.5��A�Y� �9�����w?O��(��`�����%��l��r�l��s�8�R�-��<��PT���fc�6�^>��[/��چk�҃�v�`q�|���o/�����k֥�U���O,sBg�+�B�1f8��v^ze�<>�z�����H�8�O���K��q��X��gQL}k��	����9�O<K�x�u�K �:�[�I*�y8��0֨=DX4���K��{���?iK#�Si4��I�@)�]mU��q-���]����$Jp��׃�s�4�'�����RI�ᯑ��W�Sj1��ۺ�xDX`�O4m�ˀ4{>x;]'�ZJ �>���������"��۝�7dɡ���F�!��`�pN�V��E͉�����H�[����%�#8���.��^픾3�-�
Y�7�A��`�Ѕ��Y3cGc�ϧ���u�4x���3�U3��� ��l�(v��5��: �v��J�����ׅ����4�Sm&F}z@�7�|���M���[뀜����p]���Y�W�E��T@j^D/�A#yvX�������]�F�&��*�->�@ޯ���Z�d�>%�C��A������%K���T�1y����eg �KW�2?���|[c=��YJp�B n�k�^�<_�bY�b�]Z����Rz~:0X�r����I0N1/|�5s��\�;�T��+ ���',�mw��_��T)�
{.Vd.���#����G�7��'��U4�2}F����nyH� �D��t�O�Ij��k���7�	��|tT�C/����G������QJ3�g��{��]@>�^� �$�O��	o;��<�0R�q��'L���gj�U��K�n�5��ܐ�ى�G�1h����3���S����j~���_\|�qm�
JQrXJ�m?�Y~휤uԍ��ֈ�w<�N����q��vɦ J�cjQ�o�ciң�w�~[y�]���}G����r�v��
�/r���n�t� ,)˓aʝ�2Ѿ�~��!�=��J��`M�O���xlQ�*@�����"+���K�^6��ٓ��i	.��m��մ�tMz[�߇�Pa��m&�e�}���}�"'_k�����T�L!����`����]� A�����%��Z�<>K�O9��.r�t�j1�+쎎6�,���|gԴalU�(�'ٌ�p��`�k;W6ӽ�C��q ����N�A2*��(�:[���t~��Nq��Q�ӧy��O������~^�[�v|�@��$n��N�Xd�vvW�d\9f/&�N��M/�Y+,��px�a�q���8'��-I��~#����`�7�����_S�=�,c��]T�W+���jޜj�o�a�B�k|6�k��]ڕ����Zބ�P�����:K�p�L(:�r��4,����C��:�2nZ��П���q�c�r�ƽӒ8~�ߔ��|���0�s��u���T&�'@�W�k��_l~�)3��p�O`�� �����ZA�� ��%Q~N���z�܏�b*���q� ?%�#H�ߟ�ؕV	߆�F;�%��!R[/t�i��T��^�;B��X<�Wm?	)�<I�@Ew0�w�>�1�o��0bs=�ޚ+�k���������a����!��8�ud��q[���v��Y����Z"�r��Y:�
��~��͏���2�@p���ߟN��:�'�W`)�Q�.y���{�=Y�p��o^�:�]1����ӂf"
R��6�6��.f��v��G[�0Q{�N'fr"R,-��s���IN�n��+{s]�	7�q����\Q��4�g4���Q��äX�����;f��搩��Nd��ك��Ҕ~��f�+'�	�����f:[O�)I^��=�>^�':ې7;�li��n��25d�X��h�^ɀc��7�yUe ��sU�>��������b��=�Z�D{W$4FT/n���t���ţ��c��v���|5���S��L_�x��5v�������|�%�HTr� 񌫎�s�,O�Y;��R4Ua��S�p4���_���øx&����N��45���b���Ig܂��� {���������4��#��w�,����Dz��r �9���C��ƽ��]:�g�Z5���6B���6���s��G�����X*�&� 3�;��W��Iv?�sط-��x����v��ה6J�I D�s���|W�~x`�	J���݌��i�-���V<Ałb�[�Z�ۿ�r;vk�@���(���҈�H��?��q5���/�e���SX�s,SQ���V�mI���H5�pE��;Ir�����yP0}�c,�64]��35x�H�F� )McS�*E�ʙ�	�C�+�j�+�˙!��f��0�?��>�#��s˘T��������,�ي�@h�W�V��y�U��M��g�iw�^��t�-T��oP`#u��46��g;��a�c:��Y�����#�-����;��k�����F�����3=cd�uŤ�N�nr��H��ߪY���΀�,ȅ)�X��D%Y%g�� N>�5�,�T���d�X�$FQ��%1�H��,l��SP>S���l��W�����VK�D�5�٦`��j�|��	������D��R�k��M�6)i���ρ�)bp�$�g<�"�k�S���=�ԅ��Y�&;z7���䤶$������",��1�1׃���%F����0�?�,���ˇ);h�|�e��Η�v�qU�Br8C��u5`8�1284s��w'R�5|�������X�U�hXL���0��T�R̊iQݏo�Jm�9
�"����v���|�n�"Hi�h���"��� ���m����3���%�V#�4��j�-���f<���-c O7`m���@^6��}�,Qx����36oq���,'mO#_�MZO)���;�.�Ef��t�8x�sj�#y=V�e�uFl��=�i���K4b�)&LG���S�=G�5R���zd����L��� XW�A�ً��ta�]<��;cNXSH;��3���p�O�Uf�ޘzu�-N���H�G:���H���'�<��J�L?�*�l@���|mtIWk�5}+���s3�]I�a��]B3�%�}��S�0���_R^���-1���
��O�|'&} �7�Q�g�37��oY�?y��2�7�L��A˹4І��^?�m�%TxDׂ���sFZO}K��W��ə��m� ���:Y	7��;F�岭��p{�lC���RN������@BV�eU��@*�W�r�D��
�zJ�?za�xD]�*�^������8��:�)����/�]�P��FnQX���G���`�|�oo�i\���U��� 	v�~kW��U|������](S}��y�%�=�R�s*Y�t]����Rl*�<��˘����k�k4@�Ԋ��9��	!H�]��>��Y舵��Ѕ�݁$M��� -�n�x���Ύ�c�ʺ��۬�������(?�� Z�,���UMj����A�.��'�8"��(���sК�V���f��y�X��Nc���mZ*�>}k�
�`m�iD��q�g�����S2f��tlj�X���v����T�'Ɇ�Pȟ6��Z�?�l}PS��^DTD��tA�tE��NDJ�K�E�
H	���"B�Az	������w����?����}w�}��}ߜ�2���~�n̗y�܄��O�������Nc��y�966�W
�k3#��.2��>]y��^�<r8 ��܆��(A�p���S�����;�g�4m��a%1���W����C��UX��+�rA���F7v��a�t��Ԋ y�oϮj�8�\s��΅4_a���/��d�vlVy��Z+����Ƈ�f7e�6N���U7�d���-U���R��cE-�!�q���B�z��ix�xP'�ဎp�}�&W;�8ɌD߶���dz=�ݮ[�4?V�F�RѬ�3�_�=�'Q���n1�I���^��8Z�D���m?9f+���<r���븮����U;��\�](�q����@T�����DH
Si���>W���.�S������|�y�5Y���9W���U��I��j����nO���6("L�z��������Y�㍘Q,�(`�-�#`64�+=��q
�m�zW"y�<DOW�uy�簡qǵ��W/vTVm6�{�R��J�u+=���J���[H���%�خ��?�~Mʋ�ݧar���B�Q]�zqwn�/t`����s��/�u�v��p�|J(�*z3U�*e�`b��(ҏ:�s�XW�^r'��l��֕p�l���i{��aj_>@�P��^F{�;$���ԔH�۞ސ�q�.�^���=����V�F���,Дc}/�c�=��դv�-y����]���׶_�ԗA| &J�w_�q��$4,<Rvd�Vep�:%*��t?\3���e�e��n���ݟ,�Xm�3�Y�>���3!0�:�(Aן�m���+�;4�S�a9��ܟ9k�U�7���,w�KJRe2�
�������͌�������Ɏ���Vm�W�M*�ҳ7�����ë7 뵴	Ѻ�p1�o����R17=��]�� �}�T����[�����/C�D���oc{h#'�,��y��⼖�q�V�4��["jR�����fG�����~c���{�l\�x��}Z��E<)˰�ofcV���7yKd�w@$��:F��)�SO��})��q�85�Th������v�r�N���5����GVW͝�L����`��1m�z��ѻ�����I=���������ɠg��7t����(��
\���� H�n-a�����1y��в��H>˥ؑ�)�+5�5P����`�}�]Z�	�[{q�+��z E{���xu�FAMt�i7�6�]�c����a��T�e�<��򣛣��y����qT�����Jfh@� x��<گE�D�M�6#Tt��E�����ͽ;��=rmr���O���|W�V��n��G��{:㇝��e�^�ʥKݾ�^�a{��W�drv��#�6ܿS�����1��u\��ӯ��P�e
t�$ ڞ�"hQN}Sq��ր�<^;�V�/g��ukP3���2��e���`R���8��U�]UX��W��qxM�`0�P���a`�T��T���z���Fs���JVQ��� �Q��G�f/�o��G��ɚ �)���'��_^k��V�f�cB"�a�B���;�0���t3� �p��yM���j�cv�R���>�s������t�׶�Ӕ�'��I�1O�n���3a)ޝj�����<�UK숎��ƭ�ژ��*_+�X4��$�S\5��n~�����]{��p�&�"K�K��NGm���+��I�M���"���F�j� eX���c�'�,�:5/��_V�U'U�߄��j�x �+r�2���P��0y:K�J���h�<��F��.��Z]q%�
\;;n��N/��Q+��鱠��}� ɬ9f�i���C���0���q��j��|NV�	�@�ߋ:�����χ�;P*�)H�f�l�S;TB-�\�׼�mTN-�����pB �������� ѭ��7����h��C��5�KI[AW��_Q�+��n���9j�5l������4���?��Ν������U�]��P��b7��ӟ���j�.�S�6˺��o�k�%�A�|�f@(|E%]�	�=M�~@�Dň����N���z�8�TU�k�b����w=�5ɺ:�P�1���!"��c�TD(��o3� /=^���l����ء���S��~��Tw�ӰU=�.!����5�LY����w����畩\�m�a���Mۼ�[
Ҟy��C�69�36�	A�oҭл���,�讐�N��w�k��J��9�������U?�zJ��Q��q7uw�A�
goWn���ׂ��p��ݦ��������(�Z;to�;a�ʩKV��B���l�҇��WQ������.u���W��1�����������CJݓ�n�uk8 �v&��~��^�	�����B��d�յ>����'���F�U|GQ�k)�9�0D��Ap�aJ*���0�d�+�L�p���9�L�Nr��@��#U�����J��Ϯ��O�Z�9��_ i� �ú���@��+�� ��w�&������Ε��oNV���tu��MN&����֐&Zg?ŏ�����n��z=sv�n[��w�l��U�?	�[�*���$��̑�Z�Tj��3"�X��O���	�5^����S!�O,O�R�]�!�rJ ��8�e�8�����O�}�w���$��=9_;�L��AE��uc�]����`��a�dI�H�;��Qz�W�j�Ӆ�d��
�X�r�}���CQ��Zr?}k�G�*����,?_�8!9�~u\���=�{��b�#¼p6LJ�n�~�t�Ȝ�UJ���JgU�H����e|���.>���T;�6�+���ά5�MQˮ�:����k��3j��B4����Ͻ�M^�~%�X��XJ�27�*�!�s�r|S��uՋl��[�y:\�{ZJV	ykq�2�1K����Ra?�hH91%Nư�g4U�ŷ�]u5�Q�~��>�����?[�a�ۦ^��k�dhs�p����ۢ�-��M
���7��C_A�Mℷ~�g-D)D[V^(b�'d��C?ܠ����˸:}�_�k��`K�;��X�+"�>������{����t�]��u�28YŪ�;��٤@��K�]�ߐi|�}v�g��{-NR�\b�,6�Z�$y2�EZ�8$Y�Z�و�N��4V�PL��*��WhBY�W���G�$��1z�G�8M!쩾��-�a5br�7�S�]Yg��A�+B'^�6�걗$:Yn�+�ӻ�$��pn� ��K�A3����繍���T��|\��fG,vB�g�HѭE1�	��N��1 :�}���c�����_o�Z�j��~� 7"o9�:�`���y���	|���_�n$�n3��}>8	�v�^�L�X�:�/��O��v�nmG��;�� V,l/�]��h�d�e���)�5!�>���J��g���9�D�������!�b�K�5��;���8�{�����c߇$�˵��.����0 �abq��s���b�m�����\�HЂrcv�V�n�H9D.�a�i���{<v�Uډ�56�E�މ�)c������uj�-B+��!��������&r�8��Y�&�~o�M>}�I�#JX<�%ɏ�?�F�ʍ�c:���������� v"C��T�M'�-�>a���v����*��&���!:�GM�ySܟ$w/q��p�6`u�0����$�ڼ�y|x��B"���E(�1rg���Kn���� lv%z��(b$�+�gz�������*��EI͋�g�	�zȼ��ެq�	�v��$��j���_�]*ڽ�ˈ]�*xU���Zs�!�y����:�x7I��oǠ��F�#`�R#�*��8dT{�B�9p�nLĦOҽC��f^P��C�D����Ta�n�w���wS��]zq�>g�qM?�nU�Lb��$]\�,�P+7p-r�*mc�V�qr�Jf�.���y�b�?Cud�����w�Z�s��;5�V���:���7�n��,j�c�w�e���[_�ؘ�"�*/��2��}��O�_��ue���tp�+O_pǿO1�A8B�$8��k���|�3n�B^Y��w{���J	)��o��.V��(HC'r��~�y�GS���Kߝy�&��7R����=�T �Q-�.uҩh�!�x�k������5.�Y�b �c����C��9�j^ɧG�~i��S��'y<M�9���"/>�"Z�zL�A��~=L�}!�WzHǁ�ς�~�� �OP5���<[����k���^�i����T-z�U )޹�����g�蔗��[�&��MOc)�mp����c�Ivi�cC�ڍT���'T<wܫ^�	SQ@S���P��`g�r�� �8H,���U��J�E�v�!#�������	۔T�P��+�*���(�_���kk��f��UB���hzW:�S�`M����V���@[�Ȳ��	@���x鈦����G"x=�l�q����%�8�"���c6�|��Z9-o���ڡ{OMZO��4	�L���	�Ƚ���ƵԶw`ѿb�w��
�@�W;K����%;�_��� �k�QNA���[R ^�J�哧zj�nA�~��������+\�a���WQk����xꌅ3)8}R�ILs���|ڡx����+�U��<9�#�lS	���Π��'�Q����x
����3~�x���Y9'�&U��A�>�N���VC�65�$�ֹ���%C��g}\�Ml��?8�TX'�f��|A�<��?O��G���;z����4C�SV>$�޴�Z��4�]���}�؛G����D	�BA�� R�a��ܓsA���NKWЄ���2mH�V���_g��um���Ĳ��Ϟ��1~o	�@�
|�N��F���P%��#l��q���	��X���ߊ�&Nk�����������)�SS`�"�'�Y^8�Ϟ���5y�������g4.�����o@����r����Q�f�\���'S�Y�YT��7�>���S�������'�`�o�I���NK��)U�s��;�y�`�@�����[��^����������Q��j�R���vI�]�<8�W��W�ݧ�_���=�,\c�1�q��:}�v���sCB�p�v�]H͡���ہWw��&9�{�i�k��¤f?�	oL��^u�»Q�n W�E2��u�����\�S����>�:����|-��]Xm�H�-�*�!줌AbS	/)?�������\�!�(}fI�(u�_.ڬv~��R)j�H��Y�d_�f�q�(<L��{�y���*V^@��,�'���e�2ﺠf�h�N���{3tk�pf�%� ����=�_�v|�S��˹	'��o7�?��/K���N�@{[Wm�}z�3��=�ҿ>���CH���M�N$�ΩY���W�J2(ϓف�MN�[o4�������iX�uqs&5_�B9��-5��'o��#���M���~]��ﰓ?������P�4 ���$���ө�Z��F�LI۠��E�PX������.��Zo��q�0��ζ,�e�^����Ճ3��>��Kq�?��/J]����;�nI��"Q���?����T�������W�@C8f�=*#������a��� !4��c�N8oE��I�x����9 Šwɰz��\!�U}���8ɄYy�����.){�yej�a�i�L�4�]�a�=�2��0���P�}y�v2FK�u���[,{9���̈́ەo� ��G�nƓ*U�ï����.SD�k�a����z�]�D�Y�X��87E7�g�R[�K�H�(u��r�]*��='JO�����mI�m+5�W4c-��h�F�9e��d^Aѣ�2�x�5��܌�e�/V!�0w�Ot�>����G�t�=�4|�N�֤b�� �����{�x�<1�=��Y_1:������u�G�f�`3Ъ!2H���I�&�� 1��֐�ת��h�z�R-�6���|p]��HV&��{��W����.���L���v�A����V��5g������bZ�M|oh��A}&Ng`T
J��Z���&���[��Pi�>�px?ql�@*b�]5�;y�M�T�-����~}�8Ģ��ȡ�ϝ������h���vL~���8$����
�]��IN��@ߍ��

I@���^]����MDef�';m/N4a��WB��QE�ZW�� f�����QT1B��Ewx��:㥛xk~�B=�eݷm�D�RP��E<:J�د��Q�ӽy�yw�Bp	�������vX렽;a�k��g/f꽲�|	��C�g\"�$�_ت��>Ceg��P��ɠ
w��;$�����>n� 9v����v�"q�EM���Z1�J�6������{�K�
,*!;a��:���2Ŋ]��tۡVb�,�
:�K��+4�52v�аqO��ۘC�Q{�ۼ�x�ٞn3�"��䬨h逥oo��g�3�W9��lhvL�}�3ҵƏ��I$;O#]�IF}u��ޥv%�p��(�u�ߑ>}��,҄���s�*���U�M⵹��{_��h�Sз�׺u�IV�E�Ďz�}'�<�,n��^7��Q-�&�`�qߪ���KKȟm�x�[,�"��`�����9���
[��n��嵁g�.�|���]�ߐgށ�N�����L��zj�����P����ӧ���E��L&!C�"G�XS�����&t�=����)|e	����w��
�{�_��r��+/�����\��nS�,k�O�4�u��]<�E4�cE%�a�%��P�66�C��Sh��[:��Dv!V��*c���1}I\������D٫ �c�����=@�������px|�d���sʞ�@c���u�s��&�~�4�.r�I��˱�%;uf����ϽǤ�2?D}�'�=�Ƶ���q"e"�~�����d�Y=��T�y�h�
�(�i?��[bq���>������3X(�vN�AV*���t�߇�x��(�u��_�ɣ��.�0=�W��Gbo*���\M�zK�����T�u�ׯ�d�u���ZW�.��Ѷ�SX��g��Yf+��t��r��f���u���{b$����A��m��&�A����s�tr85?����74�g͊�ji��#��Ch�V4�8��	�E�z��η�uT�4�m�g��rY�����4���~���`��A�;;��
�f��TuH"�#���F�@g��=��p�$e~��)!�����+il*6ʀ{����ʯl��i*�<5'$}_�?�&���F<�΢�]��h ��~�ʔG��%Y��#��I��+�R�ޚ�y��y��g�&�L�g�_O��I������'�֔1R��L���~��N�Μ{_:B4��-[����"'��U��.����6fx٢����܍&��5���rBw���ۮd�5��L�6�{wU{��ֵ�iP^~��9��{��V�G����u�ʿ�-��2<\��k]�Ї���Els|N��g=:Uڪ��k�b�r)�D�TP���5Ie�1���b[�<|3(\���.R�$�	<f����䒛7.��\}�;S:���fzgס�BZK�jd�w1�09��i7b�0���'����EN�g#D�ɋ�WQ�Q,s��*�+�����@��<�ȫ�;3}���|�h��
�[��$�x-pn<ԡ�Br�5�&8?%��>��5E���mb�|3�"�T�/_׶�|��~]��yҩr�UYB��_M�f b̰u�hQ��=�J�G�hر���ڻ�	�Ľ�:C��������J���3࿟�><�	p�:�NN>��T�dq[�!:a{W�I2u%�Z��{��8�c��VC����j����W�b�����Y�o������Ѐ�K�fU5Fʠ�&��~��G�-ƘD�f�+���\V1�-S�Y����GZ��Tc�L�Z񘯌Ij�W����r��컴��x��|jJrD7�H�P"���0d{�t��	���뿮��<6>:#�!hcg:�lӴ"!�l���`�׍/N�$�� A���w��J~d%1�<����-1V܅`�B�>�ȫ��2�7)���-����S���3m�ZlDu��fώ)����+]�_�筽�粁���⭛��K�TSy܇5�g��`�[��Un��� ��nV�ϪD6�tf���c�@�k�- b�^���{��հlY?�A��,�epw�s���WQ���}�=;5B�헛n���5<_�b�2V{�M�`ab�Ķ5̔ͼ�(��ҒY�b��6�W���t�	�!8��a��]�d��Y?$X�Ě��o~�a�eiu�����M�� ��QQ��W�o�z���t�:�^��H���s�j��ڰ�r��‪¬���ɃgyKNQZK�f��t���3�����훠f�r-�8�߼_<^�޶���֭ͪ �X��)�����ՙ���4�+�	K�����Cfݢl=瞦���:�	��=\X�E;���]c]���c�Q�|��Wηnj��7�)j�I
s)�xZ�c*.�Ӹ+g�
��&g��I��]�������
��QO������ʃ�O�:b��� ��b?fMN���9���QW;�����\KJ��Jc��L�~"�JY����ʗ�U,�k7�kϒ���xLc�B\�}�`Ӷ�a��:ɾ;���G
^�M���yl)<��Ĕ��;�ڀOŦL.9�t�M�m�/���]��.�,�0�V�^�GR|��C5V�D�
�-���P"8�S
r��{��\�D����w�/��\�2"e�v	(��h��YÂ���@��n��xB�Y"Ni� LuO߳a�-��Ѓ���ΊQf�*o7P��=��E, ���;,T25��H1�������o�І۵
r/�_��?����-Pj�ŏ�zݛ�zN��韜�˻��+&qה�C+��0\IF�T����@�0?Y�E�w�������x���]��)9~��kD%�=������㥛/�"�a�.Ԥ�REE�E�	3��tQ�|@4�@ൕj�/.���l$����b7�CV��U�}�&n}ٻ�Y�?�Də���N栾y�E�v 6鼤�3��t+]��[]c� ���-���݈�I����2:[HGK�_����f�1��:�r<�1�jӭ��2�� �g*�3/>��}Ě���"����P��M���<�@��?^6J���Qr6J��6��h�mP�؝�0vE�ɚ"�������F>XUR�jh�����%�Ϥ��]��n��,R�43�����@%C�Dz]!$ R���H�g�����TJ�ՃMd�כm[9{��*�5d�@ng�}��Ȓ�ƙ��wfX4��o��<�h;����/U^'���o>�GC	��b��ސ퐢�e�m�BO��,�\YTa�ߧ��� ���s`�����1��t��Կ�h�}eY�Q�} J��f����a��+�n,SVz�����	�A����ns)���5��X�x)A��4	���ɲ�Sқ����:���T�q�q�����X�l�'�cL�Q��~�cުɐub:�:�YD���@�	�M>����y{}�L��h��!��Z��Ħ&e�7�����u���{�П� �V�zO{Y?2GD�^�j��P���/��L�Lл1���(�Kv��+=�)su'�in抆O��&�e����
h�Ŗ_����/9[�y8L��.�Cv��Z��6�R�ݑ��fr��%F],In��Rg�<���C�l
�рK^��=�Wc}H�r`�A[+5���ҿ�猴&ƺ=�Iq�]����<9�Ѫ�b���J�-�I560�a�LP������mC���l�y�[��tJ� �Tb�	r��ܳt�
��@��y@�C��	2[�.�W5��.��uW�L�E�ǐ���1w=f��5ݧp��<�v����<�e�YeY��]7��p�G�~O�<��aiLQ�&.wx��Y�Bx 1���a���ߠ�����$��w).�E���n��5�'��Ѥ��Ay���m{�U5\R�Y���������� P����26R'B��g1�5ٚ�3h#2T��j�Y�.��>>QI6+�
%��E��P����T�\
L��i�2�p	9�������O���*�F%4�	�:�)��w�vo�~�Z�V|�{K�Z2J���K�߄��h\��Eb��_�+�S��Z��%�G�k�aa�iiMCOO�5��Mk�F�Sҿ˕taK��i�;�q�����$��dq[(����/fL���Ո�p]iϒ�ՠ��]��R
��#��OA=G��N!���%��>I�y����{�H�Qu�f�6��H���	[�a9�8&=8�?O*D���d���C��J@�rHSy����Z�X��Ե9��|9�%"�d�ޯ�!�L�'�qg���V���Rԥs�a)xyd��U�O��b���~Ȍ��4"I>| 4�dof՚��e����wl�Cß�d�K�_��M��^:9��t3μ��"���f�˭�>���MF�ɒL�w�$�9wt_�f��(�m x���J@r����>h�"��V���E-5�����B��Me�����4< ���F�%J�+�+��o��M�˗I��5f1R�/ ���c�:��@	h����r�K����
��Z����`=�YkT��pޱ9 A�!�@�:��_�x�4��f��؁P ��VRB��T�ҿ.�#y�ɔu�?&�J7ui�'Kϼ�T�z�P�O��ڮ�@|�Q`�Z9k�@�᧝Ǚ2x�6Wvͭ����
,˖mf� �a.�r���{�M�f�&1�����;w%Ō\�х�2�w�XI�Y�Ѡ�g#Wz@��ҍ�w��c�7�@d�.�����Ql�C�z�s�pH�k���2W�'���R��\��h�/��<?H�S���Y:[DU�Ī?-����|�?}愦,j偅�Lƚ<��C�-
dQw�-z�Ai��Z[ĘǨ#��څ>����u���M���*�@���[��֏r�~�~������F4�_�QBgR�e�a���_b��Wa��A��U���]�׎6Z��-D�C�4��B�؁��~�����t�s�BKZ@X��ݪ	a}�(ҫ��,��G��3��NOᏣXF���F2��Z����}�b��I�\��C���I�'���A��+&����K��2�����u w�k77��yC��!sjvO�1�H#0E�q�k��s�隴����kr�4e�+�5#9�骬L|t���F�g�%���	�Ǥ��uv�v���8��I7�r�8��w[\�K�:�,w}����X��5�/;���H���q5���{BC{�"����{��T��g��,�q�J�fl��r(������j^�3��_�自��y+f9�.����,З,�[�u:1K~7zA�sw��-�tyqDCٮ��,����7~��XC��߮���]��+��X��R��ڜ�H��{ct��}X�c�ʍ�k����;��'3	��ip� ē�Ղՙ��w����}��b�*������
#"����Lʰ;�*Y:�f�, WiU"�%�e!��ym')�g���h�p�~�.�iq���?����#󘶥z�e�Wԡ��@KL��\��%Ft|��f5l0#��f"PZ�6iz�u�bXA����f�P� "^��	B<��=�e�1#d����1�+�e@e�gi_Ŝ�7K����K��r���H�u�M�����Ӝ����0�;"d4+�����|6��p���j\���s�o�ݗF��u�)�l&G���e7���G�N|,ss��x[��2@�%��±Bv7���ᓤ��B��"�''wÌ�N"mg�]Z$�`}���K�R�.�;jY���FmK�x��Y_��R�� isBs3o��=1�%���:~�Q)g\����_so�O@�F���6�gLp�-f�l7ǧ����^����m"�hW���H�_��D���zx���QhW��8������1��0 P\�qA��#r�^����N�Q~fhe7�.M�y�z����0Gu����A������7��D�y4��R�=S�O�wh�2�~���W"�S$�G�AҜg
�-�:�y�[I���޻V}�'S�Ҙ-s�^��VX`��!�2��������YW1y*�k��k*|h�5�?&J(��tp��)�U�ߡ/�|�d�42��V�9���?>��]��*t0�S@]'f��4�>	�	A�G[�Y�$��sp�<t}�7�'�-6eq[�,�0z�Q5֠�.�;g_����J����4-oI�h��!�G�}���a����`N�X�������gPb�m8#�L��̧��?R�f����p��U�z�i��FO]0��BΙ�тТ�2����7I/�5��%}A�y��`G�����]w����Ɓ?��\�_��Tʾ��v�u����n��B7�	6�2P�-=xq����u���z��0�G�<�������~ѐ,s2��^�Ru��=����nK�k����N��gn���*ع����@�b�.���������DJ���K��vwK=W�(��i������Mo-�(��:��|�#�t�~u'�Sj���e��|��kCd���I&�l�ݢ^��<��z�X!���n ����Ud'�q,��ʩ�K����;Ȱ����5q�M�<2�5#���q������@�)ya~g������/}�� ��o����f5��[z�
�'���ϼ���f�[?���������o�c����K?�XX��j��4���y^}�(���;�@!���R��ތͥk��H�|�q[�|V����PYG�j�P��{/}�:�dJܾ��,pu��2����)&Θ$쩅��5r�V���j��ߠ�O�X�pB��7���%`W�p�����OC���5��gU�k�.�Sl��J���i�6��eY#�d�קI��������Ė�F���i�����,�����jr�I��i��M_KxF��{�^LįeoQ��*ݹ�l��,����
�����(�K�A���h<h���|�sj2�T����J-�Ƚ2�	������K��]���� *�:��߸ֳ1/� cU�����:���G��������Ew��Y3Z�����,��2����VVC'�t����IKĴ/ꍋˢR�C�u��2�71�l�׃ĪR�qf����G���͙�O���=(�ͼ�>@���w-��"�c�u�4x��t$��0S���uod�Bk��C��#�oAr׽A�*����3n70�e�˂�5�&)��fXc?� ~u�iܙ�SZV���oz�N����q�߂���h����W;ӑ����,�+�i5�K�"F>��x��n��R2��_(6?��E$�t�$�?s;�P��-Q"��
��*�Z�#����h�@^1��9ܧP�f61��&�~��o�}�·y�h<���)�J ��|�
��<��=Id���T�� �k�C�<yq����V_R`'=Vz#Ѡ�Jby���k��ýy��J7���CO�%\26^║I&N��;���v�8B�?�jY�9a~����F:���Bx:_����}�fĸd�ȟ&�c��wĵ\ț��s�k��`
T�e�ｓ���g7����͝
���u�N7q!�1���t��f���6�y�-z�2�N`Nk�, #����yJZ���d���W�2�&�@�:�hi���ᑭ��&3��7'K�����'�G�3aA?p@��q����i�:7�'�ȴ@��q�,6\ �m��-��:�E5����u�z�Ie�ڢTd(���;t���o}O���g��s�<��[�����ok�Ɍ��M�ʳ� 4GA4���E�Uە��ߟL�R(�됭���fL������z��N|T�{0b.�'����C����ү�q�E�}�cS���6�I�<��6��.�"*��r�x�\��/HL������0���������e�Dޅ@�&bl?Q �D�������@��O�L�g�Y��K�z}�+�.c2K�4��F1y��/�+!����o�D
�X�!�P��z�bJiO�!�&��&g����T������̟�&��-�q�h�	ݠ����j�ĉGK���ף�A�t�ϔ�^����;=�]
/w@��}���Օ��޵����P7��5�8�˅$g�N�h�p�G�.D��	������D�P�>��i��b�긭��L�2��;�J�b����P����?F7ìS=�٣�W�Tp�I�z��ړ��4zv�-���21(��~�Y�p`���4{
�V �V�<�����aV�?�y6�P�*�"$|�sE�m�2��0�78�7ų���_��#`��Jή�,�-(����=3Y�䥲Y��j��O�M�R(��"���/�c�坺8eE@L��Uڿ:�'CU�x��չJ��y<�Ǹ~f�8�ul�Lvx��E@�����'��O�l�_�����8�;�=8A$4|n<���"�@�;��|��3/R@��Bw��3Ě����L�6x �$�]�����X��}g������»�8���㙩鷯��+N5�:�Np��	�;t%�-�/?H7��i�W��Z��H�����c�c��#�)�Ⱥ���a�+�E�����p��@���Z�����(���t�N�n>��Y��S7�4u�`�TV�7��� ���_$�՟��fL�*|�"��ֿ�Җ�Z�T�������?Ś�f����i��(��PU5'A:#����'t�7����;�L髱�M�2�uJU��ܝq8� ���U�͚��q�E^��Jէ� �/�����C�,�2�;�0��X��Z�,&Y�6�� ������4����9`ҹ&���=���v��'���|	������f�]�xg�6d}&������]�s���l6�ڪ�G=�|C�¹����ڬh��f7Jh�PO�9�ػ��L�KXR5����G/<�>�94����{+�.V�8��V����߯���{q=����Zueoo�$�v�h]����b���	E��]MЎ0��3~��\���������7��<��}�����FG��2��F�j{����T�}�fJ��c��籲���rSօ�4�F[�]� ��:^X�Ӓ7և֎���ʵ�w���b��r%�^Vk�[t�O��F�{|��'��6j���u���y矿Rg�	�I�3��`��~���5u(P���.���;������?�?x>����:mc=R�Q�e@��mpġ
e����f�'�hRn�<[%�FQx`U�ɩV��R�뽗�&O�%�4�[g;��^���)d��3F����*�+���,9���v����	���G���Y]0g�j���8�d~����F����������Ҋh�>��}��f[g���<J��0u=���O�|g�F�������w��̺��q�G튄�e�|c[�Yx���e���� ��3r����L���#�Þ@��ЅZ�?�U熫��Pi7Y���i�i
� O8QMF/��[����=�w4rX��~�A�J	}6h�gk񣡍����#]G���������G��I��� �y�W��]�u)��&)��;���Be�h�$QǠ���h2ߖL��*��/����L�p�Ef��(��Q�,�r�Y\�^�q�]]!R�w5��F��$�=�n�d�����&@��	m����#g��t�+�^�?5�#�[�3������=�6�s��L@��eq}0��RQ�5������@$I��S�����C�PB�.���E��ė2�q�������6���E}�NE���Y
!HO�n�$N{X��`z��^=X�tR֘f�Sҿ�b�|aB�L"�W.Cd��SQ���ӛ��
��՚6������1�DE5��9�@ZtrY#v�f7e�Y���xN�ݗ�¶�rW$��8�r������Ӻ���.�T��XuU�"��9�ww��S��P���~�T�� ��g�'��ӯ�M��C)�2�G�S�u��1]��TB*+h�4��X21�S���=�Fޗ�ٯ&����(���� �J�7^�>r�*�;ڹ�u��k�n8+���fg�p�ya��� ��]�����:2�
%�=גW̶��i�~��K���h��h���kM������^���e� ��)��/����[���T
Q}fa�zKeC����i���ɧۃG7Ÿ�
��W��?�곣�i~H��υ@��-!a����v�ĦN뽂�S�v� ���&�Mq�� mUV��?�UX��g����?�`����l̋��!�w���2�A�^��h�/�,��P��Y�#�]�k�7 �����7�{�l��শ�3 T�x%p�3	0���2�����gE�����nE�"���G�%�M%:o��:��D��v�Jvߺ^��m�X�o$��2��H�
\�\�2�-a�O�09��)�}�Lp�4��M+�iB��-dt�G=��z��+��0��7���5	�A�:���ve.�UҸ����a��}�N������o�m�:��7Φ���}���~��ȨQ,/��&=z��������s��V-V���O��'D��q�c����ɳ� q}�d��U��p2�+�_8���{��`�^s̺�dm{ܶ%ڡ4������WW�E	��g������M���6ㅨ�Bu��Ҕzn�{�q�U'�f|�F��J����ǘ)�+d~�=m��#�� Z"�T2�"�'�ׯ�`<5ItRj�R�G�}�'�s��O]cs_P�0���rq���~��EZ���J���'����-ښ����r!�V
�8~��)F!�J�6Ʃ�� ���M���zo��lx�U� ��x3ӵ{������U'������گfk�Z_�oՍ	��h�;#�c�K��f��Q�PM�����RI��F@�EJ�D�ADJ��K@I	�n-��%'Lr�Fm���������Y=�9�u���z��;v;�����ϕL+ߋM��f$�}������+�=��l9t*����w��F�ɼT�l6V7����^7�(U7��s�/���+6�ӷ���a%�нf*���ȯ�??�]����|��s=��u2����)�	�Z�"j�:ju�f�
�g
@��Mnt'2zg�6�x�M�KN�p?4��n�e��:�b9E���E��_����gk��hK��'�u_��%���T�War���IfB�}b'"p=B��sv��+������N�|欈����>=��|m��"��Z��a?��ud�ǐs]�������.��S`>��`�[ �o��zS �I�w�R84t��*����5�U��k�,�2�B�p���]\�ㆸ��a/��|�Af1[�*��d.�$�]C��5� ��Ŧ�@P���l|�qڣ{��]i��-�kd�r:��V��mLʄ��L��-�$����3�/�Aŋ���f��$��B_��W���1�"�Y1.d�VeS��,�2p��S�����{�Z�A�m?{��Ѹ�>40[m��s&�"3����M�ϒ=[Gy��3�����v�O�R��>WVp�dW�:���**�{tSV��XMm-yF����c��%�"�`��4�J�S$U*.��1�7)�(�*��Cn,P�ao2�	�1�ު�����T�N����Ą��0^b��������rT\�Z]o��b�v�ZqIT�,����?�:�,��h��o�Cyv�M�
]��jQ1m4�ƜH�x�'�	�]F݋���K�T�Fӓ9F�f�$����Tb�*|f�d(�Њ>�3���#�B�,T����dO���w�'X�\�p�������q"7R O8�0k',Jg��玃���]���T�7}Ҽu�rl�c&���:U0P��ܦ0�aR�D�ξ�n��C_M�A%Cw�����V$������_�#�}�T\
R9�1��^tD��m��m�����=��vC�~W3�<~��M68�~�p���4���]��zoZ�$��~��v�D��&>`Uu@�^ �R���'�J�'jv4=<���Vc�r>��/PB*4�-E��Z�Q�]��w�k#ʢ�Z��c>��H�ң�-W��*�0�=w�������s�4֎��F���y/M�5���P巓�V�ڶ��i��=���&o��jR�L̀����`!�_�֌�RM��QO��Ö�[V&;�653
�������驘3M*���ԍ���O,���G#�/��
�ØK�fየBz�/t��ն�x�&2��9��Re�h��+b�L�h��>&M A�#K����n��\I�y>��e�*��b"-v�!��'�`����I�5�o���v�ME�rQɕ*�õ9p�����]�|��!�_����|E��{���Q���i#�H]p����L� {�ʺ*m6��CXᗍ�u����H�!A霮���~��&]�.���da(�\�4.H�m�' �����-���٣�)m R_-��R�H�l�ܳ>!��:r�n�yē��8���jb:�o�����������(؜�w1x}��s�5w���O~Ձ;E�LӮ�A�	vӖe�#\���\b�g�����Z�B�BH==�z�Ms��޵��>���	��}�l���ʲ�'#+/dv�`�fgG?��~��\�F�.5��J�3|*1���t����	d:;)�+.�mMm�;�/K����=���{v��*3sT�CsQB-�w���q�g���2Iz�%z���j�f��Y1�u/�� ��$��.�_��86�X�{��.�fΕ3;�֦��	`[s�̋�Vx?�)t{����8�����Z��ڃ�h��~�:92���@���@�����շڪ�Wm��6�g�%2-o�iN�[emr8s�EZ��[��z�|'�0�]�jk�\AZ��6K_�]���Pl	6���R��R}[d-��<��2V}���ųF츠S*��]jw����[wO�8��7�A����&�f�x����OO�3�#t�&��~�S�^s;���Ҫz||t������Y����
�e*����6t[�J�����,$�Z�L����m}�bl�Ja�`+��e��c�+�Y#/i�Ϩ���Ȯ����,H���76I�����zZ�|/��ǋ�_z��uB���_�"�wH�~6�ӱ�����C��uD� ���w�篚�y�'`�/K�����UHr�l�%�]����ICC�]7�S|��`|������Z�5�������G�ϳ)5S^K���tQ�����%PO����'��V��ԭ<5M���c��Ϝ��ɫw���B�o6C\�%jqȚ��}r�BLYE��չ�PF�� �ƲM�r�~�u/����x�3��P��f3��������@[���B�,�"�=y�/��	(��7�i����� ��1v��d ������%y��9Tc�?�o��\ʀ���x��z-&���,:�t<U���t��g��� E,�	�V�!+Qѳ!��S�H��|� Y�ݏF�2���y����=O�u�������u�'g��Ik���B��'��'��4���O�Ȯ��&��"����ֺ%\�2(��G`���nQ'9w����O����C�N���.�Ϯl]�0���&Q��kwl�ޝ�VT�%�˺�!'Q
h=�T��f�#}4�t���G�u+7x���P6�
�&#eZL�=-��|t����r��!J�rm`%<�{�!�Z3yalA(-V�t��c�#*�|�Gx:����zi:e���a^���Rgw��)U|�8HX�"֞{������
 "h���������=��R�RV�����#�M#Z��ڧ���^XP-�U�(��dΊ!�p������=��^{�3��.��77oq� 
���[�m��c��8��:�#�L2~��\��:��%\��>-��1���Y��p�Iq���Dt�FYU�~W�!�c@�)h�2þ���R8(ڜo�i�Y���\��fǸ�w��d�=��`�<M%~j��(�|��9��YT�Q�<)9^�����:l�������>��ܸÿZK1�/�MD�n����-�<�FC5]��u�g��-pz��ѩ�@����F��{��-p0�����E���5&�n`<>�[r-�/��&���ı*f}/��%X����q�<4��EŶ����,����,	^-���� 4�k�*��ة)���1�~�a���5�M-9���r�(�������q�҂�ը�S��z?i���������JS�?��~��4�iӊ��s��<(ziB�n_��p4ޅ y�Ϥ<W�L�wm��O�I��bҾDXOM�Bі)�7ώ1�77N��BC�ը����;q��QU�u/���]cOW6�,a���߉W/�����K0d(��hb�(}pw��Ëc��
��x��O~���R��ݹNR~�pM��Qw�OA�_Ofb҅��^��0��1�%�!���K�����L;��8����D9�-@!{oꉻ���̤r�p�%��m�)��-�um��:���U�C��;�QsW�I^5�P�������x	�D�����Oo��y�[y��|M`7{ZX�aǝJ��'ys�逸�ycCO5%�
�'gk��U�F�[#�tx���i�5C��������z�#jcׂ'�u�G��B�޿Q�H&�����蝖Hp��s��w�Ns
<W�,��%���d��ޣ�GEw��ڮ���%EY�Z|��C�^���Z����@�J�_b�KtEE��It��7Wx]iZzu"=�-�v~����u�ZQ�����J��u@7;bر�e-H�m�����'w:�%�B�G`ka�Q�sH�Y�W���?a�A��^��٫t�/��"�c!�qT���o�����ы�*�*v��(�T·����ד�&M�+�چt?ר�+膒4��*����&95�
�;YvV���L���Ƅ
�1�|���{��\/I0����s��yވ�i
|O�v&.Е�*�ܛ4)�'w?�h��y��8}��x{�OS�y�N�K�O**���d]��w���&�>�]-�Ж��a�B!��uk]'�\8=gC�<�5�yN	{/���&J��ʵ�
�U�΃� G�Y\�Ш�'�G�=�1�}lbn$�_�Y�0��H����w	�Ou�X�+�@�(�ԃP�ݭ	��e|Ry[��j)<�Y��g�敩ԵN��">0d����3�d��t >)�g�����R���>�^N��b���׬S�M��@����*>Td'86�s��j�t�%n���xN��k����}�:N���*���Q0��Z��
��Y��������#���ʢ7�?��6��I�M���0�?)��߬FߵPy�F*>��w��7�ğ�%��T�3ߍ��0����k�w�u� ��8Qkc��GX�uB2F�Q���W�(h���zx�{���C�;�4ծ	�H�o�eʞ�y���㷍y]{{�  �)���h�a���뗾�	[S�+!�6��(�@$���W�L&�i�b[�NlYkǇ ߍ�Z�K�����'?H�k{���0�:Y������6T{������N, ��M�4�^T�=ky��̌���}��[� S�;�h���]N�Hhm>���O��o�������ڬ�F�p��!�s�a�=�|�5u��Wt]@���}���� ��\��v��|��5��T��^
�9��qMu�
3˼��vt�uOmϊ��VV����9���e����d5߹
~�"N�e�s�P������S1��V�i�bO�k��>�������3\T��_�]T|�*v9�Uz*���b`�G'�{�}�<
��q�L���ڧ_e2	��WK�]S30����Se�٭5���VՠB�����A����+���4�"�U�.��P��3��T��0�a�NP@��U�7?W�K�On�>�ͮ�k1� ���1�Ą�h�4 i�m�W+�тR��T8�;,�D��
7�ޞ��0�(p�3�F�Mr�ך��'��|!V�(dVm1�ǫ1��g\�${gLP'<j���Z�Fg8��*�� �2]]N��lI��AMA��lL;?��*���a*��F�8o���[�~���JVV0�A�=�9Z}3�(0�'$J���Z�(���&vЭ��X0� k�5<OMxo����{�:�T�����^���/�*�A����j��s���eb�s�g���ُ0�������;i�]-:˳�w���>����G�~s����nW�"Y�Ī�w)K��[�j��QQ�5�H����Q� 2�谌�hzWb&�&��	�bQ4%R�s���v��*��f�ѩ����B�>;��<E ��YF��c��FN��ҧ�n��b��ʡ�st����h�HI�n'����$�3���pP@4L8��H���M����mO������2[��G<�oTw����;�ٝerU%\|:v�פ�j?>�,A2�M#�d#�6�؛K4��d Y,H\�&���\؋�FV�>�!'�ɏby���c�3=��lI�5_������#��.QB�<��0D�}t[�*�2e����;n�w�B��^u�=�����jF���|��K)W�d��.!���F�F��*J�l���x�ͫʲ�Gy��ɤ艆[��h�澦B{����M".I�󗼻�F �����'0>u-_���#����HE��UA�*},Y6�z��n��,�&���%{�*\���.�+�3�3j��M�ޙH��~皬�mf>9�6������/��9��K�3�\��@!�����FU�k���U|�u���2�|\�+���Lˀ�۠�fٸ�C��=
�\}f2G�{��P���X�rX�6�p1�L�+\I&WIf:*���Yu,��Q1�N{(�rE�)"#��e��~L�t���_�3���� ���}���e�gD���W�̽�Z)��#��o��݀(��ߡ&*�2�[h�1D8�w먀���?2MÊ�\��	��\��z�jI��؋X�Z]�XWU��ۂ��b6v�y������	B����w�4&�،��H�O�x��Q�,�z��_�����"���~�Uy��v�Bx�k�9�(�٧�.��9qP�+=�˧&�;<��|m9՘�]����K��ei)����GE��u���t���^�v9�Sƃ��+R�{��e��%,|BIk�4n��(�x�m8A�,-9�7:�&:.�@�L��09��F��[�U�>�9�wE{��I]�}okzll�H�R�)��]_waok
�AX#����R#����u�ɩ����o��n}�h�}�����~�D��:s����BK�s.���73��yF3��� :I� ��+���SJ�F�
�e-f��?�A�H�[J��������U����̋g�ʪCWK��D�f�:�d���"��h�G��/.3�]���y��8}�%+sko>�n;�u�Q��W@�&z�yU��1�zq��蜽�*���d���cJ�+�I�wi�#Ъ�^�i�_�ҵ+
�U?ƾNF�� i Ni�i���y�g�k�Ӵ�賜���-�M������d�����1,�0�[A�H��5����I���)�O �9ǲ�Yet��	4�������)rX�IJ*�f����U�o¯��;��C�h�P�Qm���|�p���L]D�>�D��K����躌L��k����&Z����<�xW�*�
r~��^X�7Q��c���g&c�H�c��]�D�x�~F�b5m��U�j�O�x�=����h�ucK�����pK���?iį�� wc_,x�[ܭ�F�����H^!�}k������M��� �]�a�4�jd�����GQ�*(m�{Cο�V��;;[±句��e�������f��黡j�/{? /��6 ��L��P(��1�Yڣc�@��U�¿jܭE������˖k���aY\^dO�R���5�x��n�4I��Sft�`5:��N�ت�&O�O���F�6^p�˴袆�����v?����G��+_BB�;;�_�)Z�8�,�����ؖ��-���4<��[����v����У�k�%����@�[6-�a��:H��c�ʻd0���o.e���0�������� �c��	PF���m����2�Wp,��h�1�`l��e�}t��O��,�G���1܆�/�~4��w���^2	w�[�G/v�����N��q��Y�y�;����uY��f�&�Y���q�w�w:V+[�}7KI���D��U9Se�Ԉ���<�l���;�>׺N+ P=K/{$��_�>�`�ƻ�Fk��:Z�&��X�@��(Z��62�mk�-dp%��#����7�p��8��?�ub�:��f��a�dW�>b+�C��o &ź��.#7 �ۂBU�
��c��`���޷��v�lɧ2�1F0Oߟ��i�W�ޠZ����1�|��F�m�~�|�����b����*��0��kIum�n�����]�:�$yeXqe;U��X���9|��V���.�}6����i~�ż�d�z�=�����*{s�0�(*�l�f�hsU\7$%�Tqz��Z�݉��H��C�4�������Q�{gv�]v.k��hu9U,�zq��YF@p�wqE
���@�e��N�3+ڜ�o8Ֆrgg87�����cMP�Q1@C�,��砷
_��JK�r;��,mB�7�T
���9�Zx]czTF��8j$=*'$��}�nU<� ��?'��TT���a���N��f@ӯ�`�G����zي[�|��ixԪ�$h��/Ο���m/�_hVy��x�O�#on�����@L��s�rk�[��q��Co+�a��%L�p-Mn*��l�T��F?2��z�������*�!I��|��SΑ;��Ԃ�Ȥ%��_d���J��[ܾsl��yު7j���������c�SX�T�_�K��m5>�k�SWdk1DGrӼwrp�+)��tI���l����O ��ϲ+~ �0�,�����$B~��]�p9� �+2�t	~᪨�dG�g�=�I��
���~x蚮/��LR�δ^i����I��k�]�Q9#m��坝RPWX@t��r���'��G��P8���c�Np��Ih��C}>SE~��.h�=i#������X��Ee�qK���<ꓙ���	
��559��l�k�w賲�0F}j��Y���3��8��q|]Cd�.z���.ZBr��sh�h��>�|E��wc���c���Ӻ���đ�?���i�V3������Oe���.��]h�]��}�W��Ö�x�Fe)���<Q��C�%ĳ|�d�jg&o^'�������~�-ջt,�R��`�V')]�tI+�Y�XU�!���,����L �����>&Ԑs�MD�;�F��ta����I�2��R�H�V��71/�D�l������=m�vy�
�t�vm�t�[�\���8�|�&������k>�i��F9cS3AA.>�C�N��k�)��O�N��Q��˃�7[� ���⼸r��jy��;7@�n���ۮ��&�V	�U*���lI�²�\΢��j{�k�d�Y�G�l���E����-"dn�eԱ�9��`E w��L�5��B�ٳ۝"����e�@۝�GI�ְ�4�*�;���n��0�0O	�%z�>��&�����B�۪��買��q��U����N�10 ���~t�K"�*dBK�;N���
��PN\h-͆lf�q�\����_ˠ�:ʜ�M$Ĉ���'���W��0I��q�T�&<P�&'5��Ej��$2��ͮ��]�t��)R��Y����-?�tUH|�E�@���x�=
�V��KV8F��ɽ��88�Mw�?/���o�Z���u�G�!k�{�C�ϸ%��Q�D�_^�L����BͿ�j6��d�I,J*�ӻ�R/K�UT_8^�=L�c�6�mli����XF����,*�%�i��$��Q8Ϛv�Y�|͔k�vy�~^u��'n�2ޚY�kUW���~���\`�RDK�U�$�v���_�揷�W�:!@�~�%*�V��eX���"^��0��Qw[�F5�	���,�7.��l�E�M�.�+쟞uY����@�Ϭ�΂��fS.c2��fRϩ�7C��3���&�u�����w���Fɷ��p�<�\��ŏ;l�C��f/�8��̠0�q��ty�9������_G�.��g�ݵ{�L��So���i��mE�Xr=�*�a_��ą�LN���|{�~���Ryh�����G ���,��g�����0�����ߍ��C��9OE�X�6����Ҫ��{�4.� O9�輸���ywPz��>��T���'��ڟ�z7\�!�Le���mƨ��H�e���u�:������/Pa%�u��Q��S�9�[��6�آD��s���m%UgZ�ܖ0���\���و\U���V�ΝJ������:�E/�-������N���앎q"�[]��2?bBG�J���L�t����"eo�����eeL��=	Z�w~ilIQT���y��E�rݪ	����W������pY8��r�����ۤ&T~�r3jѝK6+Z#u^�cз�Y���n��S�E�����p��*eq�K੯��TK���m
,[����l>��S#��� o1-
�
�^���+���{�M�˯jȴu�L��=�<Z��.t)�@���A��LeX�a~!�36�@�Ġ�0s]E<��QNK�
G�'��k ��* \�hU{+�?�a��fD���$Wl��ɩ��|�Y������d���J:(Xs���J�������fY�ۯ���*ig�$-B��g( ��E�+C�>���C���~)(����~���&.���  ��n�B��7Q��L鵫/�~����'ϊ��L�	<�`"�6E�'����g=��ey�.���
{� ��> ��|o8��Qc�/�ǯW�LtpNsb�Kx��EnA�X��	���aӅ��Օ���1��A��î�T�ޮ�EE:_�/�ªo����Y�|�ݛ�A�6a�<�y��o{��Zv+	H�S:��/�l��'��w/H������>f���G�ή�w��(�������$�VW ��6�JP��ou��-Pg�u�����������髶::�|����̼(��-d�Ɍ�"��(�0����`� ��F��XWcYD*(�d��ˬ=�s�K������tI�jή�����ƭz��"��纕�	�
�.3���X8@�����GEB�{+�K�*B�gu��Z�=���r6�땔gi����5n>�:��o�v�=v��?����L֥uh��������¯��C��m��s����G����������3����U�dGGF�-��96�)V�Ϡ��^���>���� ��K�l� P�+#�p���B��U��W�1�FK]��gJ���L�-��Lv�� ][�,v����۫Q��A?�y�_	��;�X4��Dk��Z��	�U��V���m�to�D/^��p=>͐�zpT���4������.@mu��@dY�}�T���P1�eif���q��'�s�z�ò�Ĳx[(?��KP��maæ��Z��߂����  pdw�2@~-���Ӏ�b3/�qR����c�����{�o��i����to����	j�Z�l´K"a�/���%��c�mg�XhvO,��$�<����q`|������UU��n���LV�$0.����s����jk���N�_Yz�`��F��D,G������R݋Ak��;��d>�g����s�Pl�Ztz�au�Ir�NU���+���3���+��5��KO�����?�԰�͟P�a7�90ժ�h*P>�/�H�7�2��.��>���I�z���h����Tyr�|�z7Kk�NyYPP���r]��o,�T�a�,\�2yC�q?�����s���n�%�� V��nr�"��r��$�
�d�*k��jȖe�D1s�P��.t�����B ݐӍ˒b*���$����0�0�Pq�(_�uF�6 P@�J���f�ƫ�7^��΋�$��l�Ͻ�o�K�~��`��bO�3;,�T��GS���)Jl���m.&K�)F�8Ja'=�a�1���L�Qڥƙ���:�:��ABJd��I\g�0pUǷ�D���/�� �p_�&�f�(�]�\�>�l�4e��j`��,b�	0�!\6�PZ�����|���|��yP�kf�S�#gߓ!v3c�g��gB�c3�uWx�����.#�7��3@Hq��u  h���v�z�w;�?�ΒM�_���0_�90���k����ȯ�!�� �I1B<�[�h�ii��	�ޜ�u;a��u4%P��1���]��RA�.�J��=:�̒��={7��D��ڍ"�������G�l�ښ�0���Y�%u�m����e��3; ��eD?6[���!�����\/��ǐWcݎ�:�Mج����x[T�-w�뺵5N��(�o w�i��U׎z`F�^Pu)������C�Q}���ϟ��g�/��������R�!](�xc'��l�4����9F��m��Ը�ce���zF�֙�N�ʂ?���fA�H�����i�3U�n�3H�Dl��ɖv�ZjW��Ed`���VuLN�Ć����m$e��J��e�B �(�ޣ>t?\��Ĥk�?�T� �B�F�'{XC���&l ��W��.��+�3��N��a���`��$%��O�&����+�a�;H��2��3ɅF� "" `rL�Q�G�\`$�^��M�� ���6/��.#�T,U$O1���7V-�1��,<�^�rci�����Zb�<��@�����)�P[r�fo|A�u1!��O��2�.��Q���z�$�q��Rn� ��0��y�>��M�A3�m��
^�/B/�
��מ�Il1H2�Q����WU_MuZ������� �Lz(�mk@��}�S�Dt�v	5�^�Ӧ���g�oݻ<xqU�P$z���c/g��Ő&f����������j� @�[M�Rꐎ��X7�V����z����c�AVҪͰ�x�� Y��m[�JC���]1C�R��c�g$β> v������ϡ� �[�OKYېGo}�]��҉z<��Ж�=i�t�����0���ݰ�+���P�B���a)&���S�j�<*�)
�2�~�d�� k ���Jt���!��l��r����B��Qlg�!Ǔ���W��LM�[_��G���m�r�l���Z3�W  O��}�'�F������f+���ο*�l�����Xϭ�����im#���8P�g�K����,���Gzip��0�����ą�_��u܇l��B��_�T����&�]�֜U<+
��sh��Ϡ��;`A�_��J[�xV��lLh�,u}Wb
^�閳#l&�O9�ŷ˙N��iƲڔ]�Xy�x�mLر�o����Oː3]��na�����e�g�N��Y�G�AT��V�\�]և$��j}59>Ζ4��;�^�n~q���,\I��F!�2KS��ݟx�Dm�X怿}h7=	��
�����1�/^�!t�D�z�A����a�}�=7솋d�1'�+k1�������1���On<���0�Lt��`�^��|�q��<H�њ�!� �j�%e�� ��'^���b�Ѯ�rїJ�!~+��;�|�1�-8q4xNW��;�X�v�)���n1���ԦH�u��P���:����_�f�#dqڍI�L�p�W�A$ȜƦ�t�Gk������I�+��c��Т��6�u#���	Խ�5+�H��K�`j"H��W�%s���L�<������6*��I3�}K�ی�h.]z"�F���$`��:QJ相v�Y��� r���(�<��K��7�}]�$�������/�uVVFd���-N�XlWT�;c:^�K��!�r�[k��۟�M�6�L��(��FGU���4i����P@�Ķ��.,i�ۣ��e��3����^�����l���J�h�Nx���4?Y0D�\����%�G4���T���_�h6
0�ô��g����@��٭n�L֪_t���U5�0U��3"�6�*�,�����0�y`�w�/w����їAfG�Qcڍ6YnC����6 y1�Dz �HW�u�5�N��Z��J/�@�}�^t�'�٫�M�4� �j~�o*�v�Q'�A	��ZH�`KE�I	�Y���d
O�*�DE��mĄ�D�s��˾
I�8���Z_���yi�W>2w��7�D?�^�Xoo�2���}��[p'�,`.���۟�^��c]D%6�Ƌ�;���	o�\c-�Ͽtf	��sY��]<�~Y��J��,��<s��]�2�g/���ᕜ��\:fA�J[����iܿ����2�N���/[7-�47�gl������z}��|ɪ�z���o�K`���h��р��"�Z��4/Μ\�;����7pUXɄ
g#v�y��?�P��i���v�M��jѻc�"Dd�n�:��~�8�t�����v���8�yS���ߎ��J��V+���6�큗�q+����$�X !?O��(_��]�_�>%_�ޫ^:�A���I���Y����JM�R��w�
7Z�k	�F���v��n��{h��f�Ws#����T��F0ID]Q~Ƥڗ���a���5;$���FƬE��
�i�e�q;�-m�4o����W'��5�?���H��`�+oe�篧9<󞾹�*�3ǦF9�2K��މ���N�Y?��mD�*˽!z����:&N�f+�#%� ���yNL�$|P���dTS~Ǽ�: ���
RX����ҕ(���9ۃX!;WCdvk��V������]���'��.��;�kO�_�/IcI���L�<�/X��dt�%6򥬭�j[vo�=��a�&�R�Z����R3��x0r7P
9�W�猷���Kek^��i'>�	���$U���w��rF�h �\0��X6�d| �Z ����ha����=)@�"�JY��k/��? �9-mlU}e�f�����ɂ`�E�����e.�hF�zDB0�SGyH�32?����1\I��0���m@���׋���~� ����?�>$�������GmQ��=�
N�Q^������7���~�:�9gR���w��x�Mo��r���@��
r��a5�ٹ���o��X�n��q�K}�.3���γ��&)���M��nfYl�*��2�-�u-�Q;�(�Aj�P�2�?��W�Xe��Ac4�AF/QT;�BAɬ>�`Xsͤ�,mo�����l�� �x���ŗ�~�|�ܬ�J��DyT�=ZT��M`4�T��jv��[l���Bss�);&�,�I��zK��Z3���h��>��TqΔ1pG|��� �nmt7u�k��t��osG�T���5@��7���Mn�I�Y�!��ǝ��N�_z��(���T�M����0!�z�hy�C��
���"�Q˛y%u��:���Qƞ�"��S�h����o�}���E�mlz2�`�ٸ���:���l�*4�m�V:!��ٵ1*���odnF���Ղ�e�jҨm�ҚZ�����2�����V}s�n��l�(4���[���-��aB�i��V�%qg��;��~N[2L����}��<���QF�t�^E��L��6�a;���ɛ+�O��@KЖ�1�����~�H� y��&���'����"ǍSƬ�u��2���2C'�L��<:����mI��v�9���h�3MZ ����.Dj�^f�+Ե5���o�N�G�ofj�H�d��&�!�D������Fq�Xi�fX��,�r���8���+��-\ �ܴh���[�]{��G����plA w����C@�����>�e��c9���]�v[�1uB�B����cA'i���
J�
�It��r�a\r�:�:b� ���9�\X��ͬ������D����Xf2����QK�RA�책���� ���C��Ԩ�4��V��!q�U�[x-W0���ߙ�~B���nYc\�=��������a��{��ſr�1����RO�����#}�� �1\!���%���D\\9�*w�����������:��d��l[S����~�ڹ@��q����?��κ�Q�T�9�M�XOͰd�_�J�;���D����:Nن~�Gr�<����������7��g
�o�&�l���Z�`�h���j�!���;ů2t������"^� ����
��%+��%3`���蹯����}8�O�z��M?R���8���Y�{/�KZ���W�9W�5BA \��w��w�
�待;�gY��y?N(XB>\a-�W@n������v�1	M�HXV��&�?������a 51��<�6��`�l��f�$Y�*4���v$� Q"]�Ԍ�r����
�t䣞�{�����&��.�g8g�$W�4w�N/�p����ёE���<����23��~��9�2�S?�F/*�)�4���ot�A��f\�_y�`��8�ꭣ����l�gǨ�7�v���P�}x��c�t��+���y[ҰP;��U�?C��>��}��F��̆yh5�m��߽�
��iC��/7jK
�'_�T,��"��Yy����UN�����P��{�7�s±W�A%S���Hr3[�4�X:K��He�4ҪA�]ʙ*��$8�8F:$��u���ewш/~��|����3z֡h����%�%� S^S���R��������S���vZg)�_��E�DSX ���Lc�T�taV�Z�|C_����b��j�ÕC�=��Aj�]|�H���|Kk:�b�]n�(���X��а<�6?J���G�NEVM�On�^%A��b�굜�.˓ ��e	Axi�D���0�r`|#Zj;���p}�Q=FO���-�F�����YE��.�>-j�{�9y��9&\MYD��>p[��$oь*�yk������Ĭ�b�V ���xP�ة=�ך�	�]r3�oZ'#Q�M����cN���s�
x�C9�-o�.K��B�{�ڡ�b��1?I��N��!5]�鮭UTm��K��i�FS�<��J2���T�;m�q#���;���O��E������.���BGՉ���c�$�����4Q���Ԅ�@��Ոx�aZ��]Z���a#���N�Ͳ{	�{�)��QQ�5`Vޘ��6��ҡ��M�2���\�"3���E5�ut���r]X�n���(����_fU˝w�D~{=�mtL]��g
��D�d��$��&�ڭ!㺆S,￑�r=�=�]t�e�E���l�<�z�nJ1&z�˦��g=#>�>�9p�LU�m3$���m��ʴ�➭A���"$boȠs�����n$���������y���ݹ�V"@����̶����}�ױz���$VL��t��h��f���C���5���e�=�ߞ�[�r�Z%A1*�5��r�kgMcC��dm_�,�oe3�o���������{�p���oX
N5!� F�ED7z/ѻQ3jBD0��މ^� L�:D����:�39ϓs�/��ʇmf��^{��~��޹�o^��,�r���P�������=�9%��ؖ�ł�2v�J���g�`�{�oJy��Dj˼}9��t~ӳhXm֒���/���L�����ؔ<l\��I
ܒCL9Bxu�m��ſ�젛X�@��;	s���?Xs�$�id`��^��lWT�t��
ț�k�F*emS�y#Q�=[\�D+엷����|kH��M�W�ژjY��=bX9�	-3�vƌG
nw�唰��<��Xt<Ɯ�2����lt�mQ�5�C��>O���:�pǾa��^��u�6�r@�Y�iIG��F�0Ӧ�'�nE����:��R��/!�Y�Hv���2J�e���^!m�&��s�e�S�Gx�6]C�Xv+*�|)����i��~��{}�p����uļ���`3��I��cX);@�Sd�,��y���#2��e9ƁQ�%����Y[a���H�ZW�*����|��6'�
&%�b,h��I���G,م�=�~��	T���bNg�xV3J&�[bP��\?��ʓ�Ny��x�9nDg'xB��L3�� �-V b���C}a�c��*&;�G0DY0���P^���9��H1oN4m�z�X#�"�uځcl�53R�V�0�۩��[g�5�}N\����(�h��r+��}��'��K�h;�ԡ76��?���_Z#U,`q����=#�ӟN�*k�_����Uۇ7���<��٬��>��[50:� ��sm�䀘t�7"����V�����A�Z������P��{��"5rM0��H�y����^��$(C�5Ë5�:�g�����lFB��䒐��!@�����W)Jŏ�}�瓓��?�����yf:>3��M<�2N��$P��Tl�P�Q���)>)V����A.J`Mur/���1�:˶��|g��!.��꼜?5�������y-�U�=�{-�2�R�U��l���q63Z4���]���x%q������h	��m��r�˖�����R��,��`������ۓ�j�����Hno.�k����f-��̑{.U�e"�3kN���&��e ��W��V�a�1�g���5b- P��K+܄K�P2C4�������,S*��Ag[�Kp�6�IL��s�SMZ�K��q�3��f��&Z�����nr-���|�	�9�L��=�į���]省��m��I�ǲݡ��7�B�j�0��d���cng/��$�z���\U%H�.���_����&��*d�h����Β���hN{�f�\�컩[���u���ER���^�i�^�����UFy���,�)�Z�#d��/n���($�L>�|�UN���%���"�7����Bm0�A(&PmU�뾐�=���=�7��y�Y9��{�]�E��;�u\�� i�b��(_���"��<� |8���47^`qU����r�+�TX��v,8��EP�����3;%����f����i�A��ds^�3��t���u%#�.m(���q�f3��Q�>���GB��e]�u�q�z~�vq;�������IU?�*�p#����D�2��� �l���b�
�j/��w�����7P_瞰{���촩kX߄�{�-���< A��1��BK& &7a����M'��˗�z��$*J��.m9�؇DR�0��r�׾���-���)��ۜ��ɽ���~�j�@a9G������yv�E�f���Z����ȣ#;�:��Ģ��Ҡ�&�ӻk�subك��H�#�S���V�QBD�y�@���'���R�U��$�T��0�{��Q#�"�7�oIu������߂��k�/�*�̡k_c��S��]��D��a\Yq��1Ȏu;���er�͇��8�u���� ���a��Z	���M��/���tuD~�]��s�/^V���/�+=e���i� ?���}Α���`]����0"]#!�/t�.����/���_S������GI7K��=�)��P�'�K]�Lۻ���:�
�W���?S H�DȪ듃����_Y]��y���'�Ϛk���/�D{��~5�V�!7MT�����5�� �����ӌ׍���$c��e��>���m�����b�+�夽���en����!�~�I��P�'u�:-�����R3`n���A�j�d��S-��M_�����ny��%r�f�E���oԱ��o�r��;Ɓ�E4�$Ww=6ⅵ�9���gj=M-�R�B�6}�<��,�;�%Z&��z\�?41�ֱ�,%�s�E��`�|�Uj����9K*��%�.�� ���"�Ei�}�R���i]?u�ܛ�ԥ/j�=L!f��{V#���aO8ԧ��)���!��|��W�~�X�_Iru��~~W�KH2��	8�u�
��6�۱�jM��W~�0�X??�\�)�Y�r�Ɓ��l�T^}_=q.\���Bu�>�X�v���U�����v�ߎ�������tt<��c�}u��,�~�����Ӎ73"����ҩ�3;_E���Rb��j��C���>�G艳���B�(o?C�	s��aU~b���m�����������o�w}�;y<���uX�l5b��1��r��u�ϩ�
�@�L1
�	O�>v�i�S;�>7��ouo�qU�^B����!Ӕ��i�[��_/+��U[�Y[��5���A.�u����xL�}�_|��	�u?���E��Zu'k���K0���LK%�����Q��wNy��ٟ5�֋�<�O
v�8*8;��˜؈�
B�=}e$~a���fD f�|ۃ�]�8��E��|�,d��6�g���6�|���Q�ĉ;Y)>�f�*V���>|��PKQ��l:\Q��h�m�~ډ���4oG����ߟ�tֱl<~��Re��W���'�nؐ���Hs�f��қ�,8��H*)`��}�1�/���,��V�_}��V����3orKeL���E�G��	H�P>�_>M؍%���-Q7��^a��5X��qe���+� �2��nܝ �LD�\����粃����iP�[/�����f��(%�|d�pkIq���OcR�>DI���Jc)8nF��'EE��*e��J4ˁC3�L�s��5ę|-�l}�)�}��*��5bGf��$�P�LF��Uc����>�-��[��k�'��
����"3���ny�y�GI2�NQ;�>����S���NJO�������e��6x��[H�����<��6��x��g�i�|�M��!��}g2)���S�	�t� ����ٶ�>j�s�pp�y���������1EuuL�c�Ոx��Ϧ��D��y�'��b�x�_hb�[�I��HW)oe&�e^�4��E��������L��R'�^�Xy�e��њkVB���m�4�����7G�)���n=�|��=s&oR���ӊAU}��*s�ˏ����ó�;�>�C�+��<=��@p%���a����%��z;�Nʮx�@�,��J%~�wUJ��e�rX[����Cz3u�S���)dށw�DA�o<�.2��9;
�o�|+2�yk��kg:&�4�CO�s,%dEi�4Ŏm�o�}x35`�-@z�<Mq�}��*�7%}ߜ��I��ID�����R"���)���>_�%�]ޣ[��eA������U�l��,�3D����.���-���)Ju�R�N���d������w��C������32�O�B�������TL��}�b-��m�)�^ �#�e�R��'b�b݃nSH�}҄cXq��B2�kޤO�U]gyv}+��?J���T)v������Gw���˝�ߕ%b{X�;���:N�E}q�E�:B-����Ŷ�D~��S�ri�Ɖ�Q�2�����,Gui��3͈	��d�����=l��b:�L3H�������R%�%�Qޮ�� �sd���Ϣ�g2s1�P�k�Q��Y���e�]U_N��煈v]�)�[���E�4�E _Ԫ�\rC�4�D���0��E����얳g���FS�b�p2s�	�8��T��2��Y~j��WT�<��+�Ի��0x}�{��ӈ[�z��l0��ϩk�c����2�E��7�A��IUV7q�L��U�y��)D��u�m�����p�@Q�z�pm����먬��5�x?��L�s�di�"�)���2� ��0���s	/����9���q�M�N,�������jq���ݒ~ݤ�8�@*L�I'���S��t�{I�YM2eofe���5O��u�E���g���U#Mh� >S�\x��*d�]ZZ*���pSI̵᭠�?Ne�Ӟ%�d������c��%��
!ܜU�����*~D�[�s �ɝ2�k*���]�� ,�CFm�'�~��u�[MD0��Ƀ[��������Dȼx�j��
�B�0 d^U�|�)]V��bw�A�l�O2*1�I�^X�`_����%ހǢ�f���杸)�,��d[H$��;>�o��K:})c�#E{s�q7�<nTW�u�FVʚ'���_73$5�S�D���6�Vnu��Z�AZ�q�DM��#����̽��S�B���Ȯ�*��9֮2����x�D�
8!<F�sn�e���q�ݜն�qNK��l��+���p���lTUV��C��W0s�i�k�ĭ|�p`�d���X�?8HjA� �8�L�r~c�~7q����kb�;���߂�`�������hқ�Kl����f�l�2}��z����q�����-P�i��D2���x��(�T�XԨ�(�$���/d�jԘO�>?}��'�P����C�W���GbՃ��LϬYգ#)ހ}z�ŭ"﷋���S�azt�bV7���WQ4t����7Ԍ�*�!L'W	�3���q����bIT2W�R0��d���~���/�į��jvY��O������Y&�����z��/�lgs>BK��U'nR��཮.��_�>3N�+�o��<O�A�Y���tX�"V�o��m�ٍ�@��<b�*��PJ/�3_q��̋X�};��`"k����Y���Z�g����㵥�T�_���9�����Mҥ��4�A���Cɸs�ri�UFV�?����+8r$'U
�7�m����GF�Z�\��~��HhQ��3��_�RT�;e�+{fU�%�ӉAw�S���v�sGd�TV�G��[�M"	r_/�ݑ�<<=꟔v�n�i5ҧc���M;L����8]��Y�sbf64L�mh��x���@m�h�/`o��<�0��Q�i�����+��sSu`�l1�U��I����0�O���a�!���||a�`���TP�,R�j�jϸD#kH��e��K]D�g��'�w:tQ�˜\Y��̫%tFɰ�e&���J��<����	�ei	� �]e��!�!��xL�HpM���P' �Ⱦe�N�}�0��8ei0�.lbˑ�M�G(F�sy�P~��=-��M
�<�8����(���/#��:dfl��i+|a� ����ʋ��pxz<���ҕ2�J��^6�����s���0@%5���؀Oeɍї3�0��b������8��Z�0��� C���7u�M������|9�c)���ga��R�Ż��1�v��O �z�-�{�W''����˞B�:0x�&�Q��Bӆ��!�2�&�t{�7"�M��j�C�W���_���S��Rڂ��qkѾ���p`�cnH*�.�R�!���]"���v��8Dw�wn��Z�(��Щ�'��:�-	�3�Jm~�:����4�l:��e��X�]�1u��tD}��?E��I�X )`5�D��u��(�nX��ݰL�3՞�������D' �����JPr>����	���N�-#�԰}7vMy��I?�^F�#q��������#K�m��g;�B��&���G��	��סq"�Р��&�aMlQQ�	�_�j���e��]E��I�xq �d�L঻�Wn�-�����4EKFk��|�Nk��Jb�P\����0N�ю,@$m��ǡ=���-��f����M�Oq��\'�V�6xf��ᔋ��~jm�!��Αv��*A�T \��k$�tj����O��ƔŢ��L3�{o��!�Y�n�PPΌOW�U�>��:f�!E��a��2�(z95�<ŽV��@����{s�	�8b�2���;+��:�׶�0�ߴH�>�i����w.*;�!$gSd=�ә�ڍ{ʵKlm+�G��FI]���c�
��~����$]P�{�Ub)�ڈ��g�z��Β���*�95����qT�n0S���Ǯ�j]���UP26��?�Nl��	ʑ�/�oYʯJ[S�:Z*9:��?�J�*��NjK�/,��!���5H;��y?��lb^���hf�<<go�)�]�����5�]�k�0��-	�"7���V'Q
�/8"`>��R�7��
���Ą����B[��z�%�a�H��>�p�/
nH8����7!�-��&4�7L-�M�w[l���U$���(x�%Qj=V#!�Kp4��h{����h���`�ӕw/�X��4f:�@��u-�B�nEPՊMu��f�DV�7���9���uJ�{����,����'�IFG2�J׫����.��{EKvD���NF�]Q�ۯf������Ӛ|��*šAW��ݤ�ܤw�HS2�нj�dq�6_���E�ju	�s-8 ���0-98��3_�p�W,�up�2��;>݁:o�婒9MН�.�T�W��ދ�Xb�^���Mm�ud˄4��*�8��~��_�2�|`C�;�v�}^����n��*Ç�Q3<�=�:˥?��L@���>r�R��+���$[9-���r� l�1 �V�x��CeӅ%!� ^�!���9��o\Y+q���J:3��K��7]<.���3[�ZaL��$�V��|��B�MI H�!7���u�+׿�էF�h����+�d�ݪ��CGt'�}Z���KdV����X�E;u@Me�� `n��3HS��?�[�~ڬ��n�e��������_�)dD3A�
߮�s�C��\o�oTx�,(��ZʅoQ�8q�EIs[������>̫Q�����?^�K55�l'E�B�1�+�c�� A�mIX6�䬱���Xs-��Bl����� �d�jURXa��)y"��}.{nع�j�ڡdR���(l���x�VīH����%��4��T�p�^����=N.2�h+}��>h���&7�� CV���y���q~�����#Jk��t�C9�F�,���68�� p�\�����3^*�Z(/�L> ��╧�R�]%��m����n�L8oއ�K�U�13u�Îͯ]��ĽS�7���Fs�t�;��1U(=�Wi�W5Rg˷�n�8��熰f�8��Z�h�*��JN������6L���E_�7{�B�Hɨ;H�Sv�Tg��,x�&_�h(-zde�k�/W��PՖ�������\��2��`Qx�^5�� ��� �"����Tw�)ą�暓�\Z�,~��:��9xb�~#���ٌ磐�}����4��mɯ=��4�����TR{�c�ʱ��\�ڐ����������Q�O������jxVf�%`���i��X_�3��]j��������l�כ3(��]��"��! 9=vI3>�%���E�ӄ1����H+��$����B���H�Ś�M�0�z竾nɫ�3p��^}����ƺ�ҷ�vi�m}�NW��������U�i�L�=M�fw8�gd�,b�h`�A�=PR��z��xR�'�:���IB��r~���e��ݩ�$f��@[3��]$���I��L;�&r!�f�L��}51����V�̿��A������tU|gq���+�w�H�g�I��"���Y����tz��=̥��3��L~���r�qE�qQ2:IP��h)5�0_6���T@���<��˫��/�\Һ�96F�I��:�r��I�94�Vg'�c��!�����$D�ʙ��:_���0���Ȓv&�ElZ]o�5Nε��4��R�M6���T�Q:�9�%]��{x:�O%��o^-�aп�hB�DUn}�|3��Q�����ˇa#S������C�`��V�V�Ѕl{��~5�K�~�(��'��o�-A�Nj���������i�z�8��u�i�h������ҜV�~����r�T�����5���u�����&�ӯ���7�z6��g�������i�#�Ȣ�n���ܪ}RD�9�
y8v��K��\���p���nK+hJ��F;��G����^�T��"��ƌZ�B�Y��J�g �Ի�G���d7:)���ejw����N����ư�?*UY����j-vdg�+Ґ�-]e�6G������s�Tl�L�w5�Kg�a�,��94*�q�Dnמz)���ƲJ�@4a�ˎ.�͞�îFԌ��zd=wg/���/���t.)	���ޮ��/�󏒲U;S(�M=�Ҳ�:�9�̌����-�OT_;T~sb�����8(�,KL=���� Mm>n �g*�."`�J��o7�	B��Z[����z`��>�F��o���3�������v�q}����?��S�)h�����_��R���h=�5H�G�8��`�ZI����J�(�:iC�/�uz��ğJ���f� 1��V�Ieǁ�[$�Z�����̥%�)�"CY�-����Ϡ*��.�����Q~h�����WK(����'{�9w�&^D�l�`��_m>��I#��ՠ����v��M�+�q�ؖ�C��/P.m�ө�noУ7�-]~��	�R�M�q>��9w>k��O�B(jnN4�ZS%��G	F�Y<Ե�����^�f�1���&k���7pY�~k$�8�_]�?L����~o�)h�I��}�w��Nb�0�r(���2����P�T�ϒ2�X��.�6��CM��'��@Zp���O"�&�c��Z�5��+i����W��:��1�_�����m&ٶRG�2���P�:=[>h�P4���_3rdY(O��
G��PH��c`�R�LDt`_�uK�g�d�}}���L}B2�fV�e�Ō:�{+�5e#J�t���ɳ��m�n�<F��J��#�c�M����>Uk���������1U�$���%��<=�*�j<���U1��d3y�#�l�D<b�S[n=�%��̘SG�a8�rw�뿁� �Т�dŅ��Z�{�}2�E4=�"u�n����n��s�ڊc��}wr�+��֏�^��8B*�%��k�ވ�5/���A����n�x�-q�4�Ҧ,(p��x��	�N�}���ң�6��?�wC}5x����pq#,L��}�⷏_^���/;�6�6ݽ�I<Kuj��ǒ��LD���@���.~
�_J7��֥�H����c�S�|���~�BR�}��l���%���Y*3q���\�~>&%�V�b^S�?{�t��M��۟~����_o��֫u��t��Aü9�E��k$����Y|o�A��� p���[��F��M?l%ھ�ȵaSQ�!��\v��F��eݝ�
�b�"���]�R�t=y?Q���Z��5���%�e���i�_T'����A˼�����B�i:G��fQ	�L��5*!�=I��H���혐��9�ЭT��wS�^q�����?R�i �4���q�Ԡ^l!�s�\�4&�^�^E6�S�n�d8II�z,RH��Q��̴�wb6��+����PY��J���1�7Pj��	�7���Cz錛��K��/�V����[yg����ݑY���!���K�%mɫ�P���&Â#��7iX0�,��d��^m��,���˺�������qQ��U48��8ujhg�̄������_����Jd���12R���R�i "Sz�|�K��r!���	��ǃ(�a�I^��3)��4��R���јnG�(�iA�f�;H��E��u'Ȇ7�MI�4ZoK���r�0t��!i�ޔ��� �襆	�&)̞q�1��e�k�Mq@/����ݒ	�O���]�>D�4_�bS,�3�T@w3�pMϺ���X�t}QI�PT+٭+�ǯXRl1�΅O���l��G�#ې�AI�.�ǣ����.�����_��VV]�P\�i�$|\쿣(����Fؾ���/�,�XIe��d��h
a�0";�$$#nr�8u6��
T��^��^@Yax�q-5�WɹOnX�_��ҁZ��TXܡDn���ߐ��
tl�I
/�ᦕ�.iC|5�ʗ�b��l���&�5��~�כNj���������F���lp˔E�Ű0�p��n��QU��@^Y�U�z������7�>��?2��H��~{�J���ӫ�����r���|̓��ʗhL��Ť�A����*�-y�"*Q�.��|kP}�����iX���������W��-v��A���+?��K�Ӂ�E�&]qt�MBh�J�\ #(3�Wpe_k:ҏz��2e+��5�:�0&�)�>syN�i3�'���j��-
c��d����~�V��St�r��%g'&8�ށFk����t>�����hl�$�U����l9	��*Q�44��a����<#a���!/V?̿q��%[y6�0����`�G�r���rDҾ!�V�2����]);���?Ζ�1���� ǳ�*�J��/�6a��2i1���nʑ��Z��hU��DS�Z����G�ǯO:��q[|�9y�&e�/Ȏ���+���Q�O-J�������B8�ί+�0��]�zQ'ʁD���V�R�4)@��Ebօ��e�]�|�5�Fԭ���T@O�*��0�v�U��ޣ��	�g�i��TL��-(�W%F.V�Ĉ������[R�T?
��0Mg��E")�ƿ��Sa�2���\͂j����١�+Ղrp�|��Xז�f~�K�����(����V��w7b�=[s�(���[�)��Mο��|���lm�L[Hd`&�y������6N��q�����ͨ=��~<����-�^�	N����I��54�^Q-p���eQ����<�J��mL�Ȩ��6Oޘ�O�JZv�b��	ف �d��܂Lu�����xe	U
l����[��4W%r̵�H����n@�a�U��W�'3�/�+�m�X��*��}�m |V�� H21���Z�I�!����-c�ĥ��<�
�82��=Gr8�_��čb��,����or�~���ю0��=����+�>�Ҁ��n�����n����0�����vg�k7�0�i����Kɑ�<��~�(��/��خ���ctY �Pݺu��R����P�1i����n����*Gڨf�U3�7/��4cl����3{J�19�b�uq
0?ċV��6���	�����O��8�)KYt�pu���Е~���h�+�r}i�M�c�3������T_�^i����2ؘ����X~~{��p��ٗNE�W���k���Z�Ǵlt�Z���V�F���_��l}�{2Ԑ^�&�q?s��co���XTJ+���ȗ�J���s#]��S���b@4zT#��Bj���5\㗂ܺF�>9�H%���r{�M�����QG�Y�U�O�nqs�-��)�O�sl~������:�T\H�����y�H�(ҳ8�q��f2�S��H���3�3� ʫ���O�mJp��'h�:�t�xv.�nʿ��E9*o�}J<���\ϋ�������#���TE���q~r���Y*��T2�Yc�X �=&`qh%���p�g|0x�i�~qA�.�zh���o���Wu��4��1����5Wx�=��@
v���DobS��-!�]�+�8x8Xۥ�	�Xu;<z����:�E����̌��0��Q�fwץ�T+�)���}���x6���#���[�����:�b�揑��tY���q�%��-���87B�E���L��h�D�����n
X�]�0շwL��˙�o��B6q�!�a�z����՞��9�Uh�C��+��z�����ЩP�=����f�%Fp����$���R������7����+E�n��f{OJ��vsW�-4�n�N�}|Q/&ӾI������u�k���k:�=��#8��X���>rh�^���rY�F��f�J�1��?F:e�r׼ji�.餩]�|��jDL�Ejw���W���˂�um�$�2�M��0(���������΀N�R7Oʠ�f��/��.��6W�n����Cy�BNEcj�Z�p	���P� ���?�c-T�]B.����YZy2�3D�6͸��ò4Z#}W�?�]H���A���sy������c���RA9FM���LG�?��n��\���x-�U��0���.���ދMOj�R�9DV^��Qۭ*�vgH�u�oBR�8o�
g�ST�����>�Ȩ;识�U����V���X�����?�� ����4����hpq.��ʓ�Hv�ݖr�������AgȾm�؊Nђ��u�'���T����3R˔��)&���	��:=gB�\'�c���S;�\�:�HQ�R�����*�-�xVO���B]����{�������u-�A�d	֦ɱ6�S�ň͢8�?�%*6O-C�@%Y0rX9]�_�Ԏ��؆Ù}����`�%��>�u�@:gI����3�OϞ��t��������zXA^��`'u}�u�w�?���ʃ����ϳ���..
��A��#��9��e��L�?��橁����M����,��M����y��Yh��&�v}]�Sk9�TK�^��x�*�:�+\>�rH��wR�?�k�n���*��B�9��l�='*��`�|;\�f�~�~@��k�x�#O�V�Hw�����n�Q��0Ƒ���!�g'P,�kU�fC\�L�T�N�(cž��n|_�c	���۟��,��e�S�:�6�6��9�����1�[�G��ٶ��p($�7�v�N�K�gbn��=Y��	�� &�p�eAb�7fEB��_��gvSd�U���>��V�b/��z�!�ĳӍ�M,�1Q63�ς���w�������!̾b��)D��眭���`�Wn[r~���	��caXP��VU��HG���Ŀ/����QX�f>��V]J�{ �\	e%O�RPs0�385�/%�F��?A�L�G�;v�pH��b��Pu�`���3g���i.���!���g<¢��]/�ӹ-ef�~�Sܠ�Y:��d'�z��9[�<���ݴ�b|:�	:8(���sQ�^|cE�K����~)���T_�;|?W�^u��Y�r>�tX��kF}�5S�9z����R7V^��x��Oڔ�h/�]�!��񨷱���Q��ѹLڹG-�e��T��S�x3����;�b�P�Q:].%����9}
�*R-I�ç~&wx.�f���}d��H6B�X��{[��A�g����)�� ��?ul�kCY��7��J���*�E�?~�)�i<�]���N�o���E��Xr�o7z�&Dk:
N��I�6�T�HCb�7L\P��K��g���E���_)H�ٓ_���e��'�f����Ik��S�_����WT�;�et;�Ӯ���� �-��k�4]�_ �zF
ζ�������p��]`5�_�0�i�)"t�H�|1gy8�7U*�6�Y�?� �?��,���0��,�)	���k��1�g�88� h��g�v�U<�-�E���۞C	�ӓ^�~����<#���u��-5,��j�JW�>@���7�GF�Q�R�����j��Ժ�m��d�g�����Mx@�p�4.�z�D�S!��_C2G��a��żv�ִ��/�"Q��b�������a�e���ӟ�i�B�zцg/<Պ_�~�X�[�	*�@O��Շ����^�!��х��N,��I��-�>�+%���W	���?��Xp�7�r�6U�P�Q�5>@�Չ�Hx��W����}�܊
���T<Y|���s/��Z;�"6�D���99rԌ�}X_��]�N_�b����d�bR%�{9��x��Gj�H�F~���=lRH��{�УQ�Tv	s�S�b��M�ӟ�Ir�˰E��O�6�&+)��q�^(�`8��ᩕ��-;�zPK�b�X:�,h�Љ���4>�v� RpHf�����<�s>	2�ߝeC�,ܬ=����Y*�a�L�~y��[����r�Ry|��}D�"M�K2<m1�n[�9(S.P�Z#B��J�j�f�2����p�sOi��1��`� �3�-�EsC�tY�a��7U�B߳5��g�L�4L"%S�#�D�(e��h�j�J!�ʴ�p:��|��TN�ߐ�Яz��ݞBE� �W�1U����F۴�'�\�ٛu��M6S�j�Y���	C�_"���������K^�jf�mH��[A�� ��z��2���O��8�7�BO���F'����ow��-h��ht�Qk��z_��O]�����(��18/c�n8��әGz����G�����޴�V�h^?�K��w�hH���:�����)6yOKT�2=��,�u�"M;��}�j��Bg�S#�1�c3q978���,G����b\��:d�;e��R�׈fN�2h7��0���D���E�����7XNy���%VQ��ޛ:p�Sִ�"]��NE�)#C����P,y�Xve��kU����Ƴ4�Rŵd��;4P��16Ì,��!y-�B��`9��u�Ln���4��m��Cgː�C�C��`��z��H�9�}��1�f�Rb���o��א2g�\��LT�Om��
)M�5���AH���B�|e��!N�.0楝�O.����[��R�aKw1JW�� �W��IYIf�煾_�.J	�[1F5[Ō��)xtk͚>0����q��B��~U<����h�B�shwM�
�q�>����^��k�ܖ�m<:B\VY��e
h?�sw�q����If�k��[�4�W6�����Yz8��V�x'P
��,���l��w��A��DLOى-$��x�t��ڮ�Y��g# �8��E�Pz���礷��ZB�(�š�hEtIn�����vy{v������,�q(�nU���9�x�B�5�{���3$�&��z�ǭ�h	{�Ʃ��6a��������^����,W��rx���]��y3c�}�7O"D����gNFc�TH�mT�ei�Y�?%�g:�T��D��fU�n���{	���I��x��Ԧ�����}�� Y�K)˨nu'��0�(�NL�ܷ���a��^��~�oݒ�q�#�_բ�l�p�W���Z�6Y�yƙ;����SK{G^�䆦��-W���_CS�l��W�G��{)�=���9�8�W2O\ɜ,R��leaf����>cm��H��WbEJN/�'��Q����L.u��cI�M�sؘJ��cd	q�:&�h�o��,�i)jL�#���WF�@�R�^��i��/[,�;��١?�ݳ�v���Y�l�J椽ă�F��ך��<�0 jā>66s�}���R9��e�q��c�g/��C��?��'U�LDR�� t�+j^�_�(�ۂZ���t�Z�١��lb��ƒ��[��H�M�8n	���d�c^��%�z�z�2KV�ʌ�v3��\����h�,���^(7��>���~�Z�������-X�R���q���yi�)��i�ꈣ��s���=��,QC <�������N����d�@88>���? ���Tՠ��~��|�ty�U�;���&eIEOѲ*t�V��d.�:�@ʲ���קE����w�K[_ tM��\�S�獣(
�Rc�G+�%X	�E!���~ ��|�[a�Z��	u7�[�ͬ�.��f����M�SM��?�;�=�0́����Fw��G��B�w���I�.԰����� +L&%��T��3�a�I���tAei���s�w�,]$�'�ѝ�b�+��Ĉ��,���M��e�5�Ҍɫ� j��P��x� ��o.*�F$ŒY�>������T5�X�_k(���ʧ��x���S�1>"��מ��ɭ�8_�\w1*̡����}����y�qfّ�����H��N�9E�᠗+�n�����vC�x�eA�u&���c�)vYq�=���(�Gg�Ӿ��l���EÁ������oM:,3���m	�	d?�pϗ�͖�#d�A��r�-�dUJh� :W����������P$�����@��U)e�C�7�X�dz.���g�d�nE������T�R]��X%0��/f]��m�j�㨴ݰ;g��;����@��8���ws_rc=��yrn?q���{���&,ψ���]��l��ur�VIxV
�n�$�ŁH���`�h<��t!J�j�DV��8uIn.fV�j�AUt��v�4�����l㈦5�������h)S
_h�j��W��ni«1�Έ�5cʫ:}��?Q.�R�uH�^���7�@G�����SLL��E$Z֬ai����F��D�eۈC��T��Q_��|^)`��xZ����&ڜ���["_qV.q�d$K1�7�m6j<�5�������x��/�3�����#q� r���3���㻋e�J�8�x��\�W�����d�HF����b�S�A-7o�.h��s;"l7Η�~V"���c���g���j��)7�O�1}�leg��-L�=�o����#�ٔ8=���-EEF-H�$�0�B.�)��J�b5c�BcF��L��IS���N4RtSI�`e��_�g����Ne��%F�F爴A�2t�٢���+5�3
�N1'���L_M1�nΏz6=���,���X7��kX"t�Vg� ��Z�䟧���0��m;m�s#}�����ｭr6�~��{'��.����D�9�-��X�o�Û�;,���_�m�f�+{}u9AL
��av7��a+̯PK� ��T������̞�a�UViV�(�R�KgD:�!@�C@ElH�^��J(J蠀�H	���K"5@(ϝ��{�����+�̙3s�53���+�ے'���~���y"�~���W��\$ڶ������x��������w�@��d>���C���$��;�PbXjl�t<���0�n��+4>�$�c�^H�6j�ڒ���&;�hS-�F���������%H�2�RQ�i��o{q�['�~�_�>!uG� !r����)-[ljh�rέ^Xo�q�:�g�����Qn;�w`d�1�}|���逵B����G�f{�Ƚ��������}�ɞ��K��'��y��&�6��B�tc׸7�{<7��<V�-������0�I�?�����X����hi#��'�7�`��N{������@~|W��l�r����j)a
"�-�,����9[�����V2��{�����4[� ?0F�'0��z�2���e&��_�݀����ZFG����N~�Br��"�Ux��/.=1QOq>X;Q\�����)�~�y1�_����sf�j��35Ʋ@��\�ʊt�..��&��\����F*���ƥ�u�E�F@���ֈ5�<"��z�3��K���k�����[�@$:�H�-X���Dń�}j��j�2ݾ��Xi���r���˧�Nn[���{qJ'�)�B�R�GX8�4�9OV�o�'�Ç]쩃�n�����eŗ��L%{��x+��MS<��ypݡ{�2�Vq��2~�Mm�q3B���A��v��dz�B��d�U��]( ���Q�wґ����P�/�LV^�;�Qys�_�	��k�1^����6�~��0�W��ajK��(F�z�"|��־�F�$T��-=PA����q��<u��Y�&Cy��Z癆E�qX��3�T�5P��J7��hI�чC�KKlE!�>Ã-/{/�&��5������̼�����~�����ΉW����S��:T<�k��]!�>*�������F��z�9���41��8��x�-�x��!�>�>}S-���{Ve��	Tu���N��G(���H	H�;q����<Df�n����U�Oԥq��yD�������e�4qt6��~>(Q�5�g��!�1�#۷YmL�^	4ۉI����O�������<�s��9J%�����҈]=����\
�S'�፾��~������U���♵�3{����T�/�~�� ��c�z4:�MF�.G�T�ѱ��щ�a]V�R]�+�8 �?v�:�z�R�#?���RC�{P�Xo/IL(���7�4=b��Հ�J3�e���y~���֩~���X�^��3���ޱ����f��o�GH��͏z]!+I�>��jC5{�6:����8�N���	��[�GһXq����=��re�߀�f����$,���e�}xu��U��,����F������P�s��X�̧6���Bb��7	-�GGQ^������$'��Y��n@�IOY0�d�<�d8�XA�W�ko��u������ʲ���[��#��,,�̌Uj{]��=�?D�4��v����L<�����o֚[S�ŧ;�U@j����b�X��P�< ǡ��Fq$�sx��*^v���YM#9k�w�w��o��+3��'�ф�,����	����&鹼�Tc�j<��^>|4DX�CK�)@ȪpuM��Ad�8`��f�����!}�����d1����X��=o�4�n4F>B�Ek��{����@�hHb�^d�	�z�AH<�C��PJ�ݮ��T��C��
����t��zUl�R0O��t�q����<��|4!en3�pJ����d���p|����2O��ń�Rs��k&c,��*iu�Y�(��ա|���څz� d�ΖY����/E������Oa��+�F�j����=�R��OT9z���Z|���7�7Z�?L�Pn�C��T9"g���������M'��c������=�3}���L���+TV*����UF�P��T�*?K����B���	+��{v�����)��^m9jd5u�8,ĸ�-�b��H�t���h��:LF	`�4쒤����	�Ĕ�v����7�'Ƹ�!_:n�;%H���o�l��U��t���}��)'�:bzu�'��;�%�=0�\�~x�;x�ܜ&�����/�l~��G�k�+ո�ܺ�&Ǫ���+��zmz�^(��$oD�=8.�� �-�^�~��Cr�{M���'�ķ((}<�@Z��n6�¥M<||`]��K�>��bx�zPEn]w9�Gby,�^��G}J���)r���"1�|����'�0�2{���2�%K�s���*�i�ٕ��(�}�zd�8��t��>��&�m�g~�~�
նZQ\�#S�F�h��ه$(�ZU��(�#�.��i���W����4Ѻ:wȌ�~,�Y�c^z��c��ő�^���K�7�u�y50��#4�>}VA�v"S#f%����ۅ؎������X�p���Mr9K�ݡ��E'�Ā�C��������(�TI.	�۽��`��5V�JU3}^�~��vY��ZG�\C�">0�9'uJ�;�o4���RFܫ`X��O5&-!/�Q�.y�>5٫�0���2�f;��.[6���U�(G2�� BV1`eYZц�~�����)���F/���h�N��:uNn�sٵ�厠��y�������#��]o_����6���e����1�#/]�����|��ջ�չ4�v���~���P�a��Ѓ&�;Q�w�)[�����O��*B���Qn���`$� ���jtU�ã<�X��Q����k�#��p�y.��w��EEH"�;m�P�k}�0Os����[4E�Ri��3V�#E��=|�����Һ�(g9i����w�p�6-�f���Cd��=�R\���ڳ�0#��NQ#�����p�s�S���o�V�!������U����*_9������b1��$�NQ�@��V	�K�u�����o�y�l$;�e���ϳ�U��ɜj!F	9�V��ݗ��.����D��/�3_��
}8�^P�XN��b �������z�bcޔJ���r~��jhvlW��7cxs�C��u��Z-�r� �����<�R����S[��y��^wD���M�[?P8���s.%��Iw�>��l�W�J���FEsN-RO6��> ��$ؙx�R�*���FU��.�. ��A1vt��.:襇8�`�۔5�T9��t��	cr�C��a�u4�G�+g���W��g��E&7��K��84��V{��;���џ�4�߲�E5ZH��FL�տ:5�$v�f $�EX�{�r���b�6��x�/w#i潋@�.yv��� r��ّ�a_	���`Us�9��������L);_���8.���=���ȠI���v
������hN�!�������g��	�M& .����Ti[ߑ�^�#s0�s��T�+�v���}i�[��/�A1�k�UI�h�QM���2�to�evr-���v/���#���Y��t�_rT7@oV���'�M��(����p3�N���|��
wD�P �1.�2(�=�c�̙�Ŕ�>��зz������J�A��ސoP�bh��Pqb���"����]W�2�ۿ�JT�i�wL�qE�1�����0���SW���Q1��3 ������;�a��ӧR��!?�u���9c}0�����r��7B�����~��Z���N��s]�c9L-���W*�ɵD�@K�Ů�k{Q���W�>G$zAH+̃�_�U�B�RP���v��#?���^S'��:��~�qEM�����E<��)��E�Ԯ�a����.��ħ��Z3W�<v���ǔ/��\ĦZ-\ ��������p��
�G}�ە�u׭��2q����Q����l���}�`����<lڙnA��g��}M�
筷4-�g?�MH��2��Q�.�Q���T�݉�;� T#����`^.��&����͒�*H۩���TC�ia�}�����3�r���L�H]�+`<�*�^G�
�[  �߉l��^�mon+��|�"��ŀ^f�)�7����l1R���7�h0QXC��u���h��zG�-�և��0r�f��˫L5{s*"ε��R�����vy��xB`X��lB.�W���;�~p�>��n����;���zM�WX� ����8F��Hߑ̩������ȒX�Բ�a��+��	6�[hW�t%@�tR��Ə�&v��Ét�	��&��:�,�M���F�� DX�MJ�&���Zۥq,}˱`1�D/��K��E咴�V#��}S;K���i�K9�&�W�1|dJ���q ��O�%�q��L��V��x����Ttq;��f�j�!-2k��*�
�dNr�iP*��Bkk��
n�}WV�b<0 ��
������i��qҿ�B ؒU����#��Ђ��UZ����:�LTg��������V`@�q~J�����X��2#Ӏ;���9o�r&\w��9���u^17h��)
�4ִ4` ~�k,�Z"�U� f�� -�/���{e~����$���T�h��8m��Ɲ�''���2�C�K���A�߬��q讶�����n*e�n��G6P��ʸ�x)F`F�I/�(,���D̠�r��r��~U�+ kX7�Z������EIZ2��W�&ҫr��ן������(�U4V�ֱ��W��̩�O�|��m$�"'� 4+��v�D�4#n��?�l��� W����X�I��;]��kS"2�˸V�E�������l�A$y��Aƛ��v8��Jw(w<���=zt�Ⳟ!�u�v��R�(�"�w��Z��L�xH�c�=�g�� 'o�I�> 0A�a��^��$��-�a�O�f��ծ�Q�G����������l�;�ĖZԾ�i5��y��S�І�9�� ��P)Q�D��cӣДҚ�S؉���sh���4Y�"{�E�Z���5��Ch���γaͭ	i�z9�zS�oX��i�c��H@U}Ҟ6�u}҂&�L�}���à/���Z���iX�P.��R�噵�$�鋁�wgg��7$��;�[���|�/�#?��.�����h�ꄱ4 ��3���,��tc���	�W�WG+��Tyt��{o�9Udo�	�H�E{pB˙R��I�C`i��6���˗2�e_O��9�TJ�P|i��~�a����ѱey��Ch��fI��CS�w�@��C�1[��=.�%�8�=���w|�z%DCcȍԷ���b�O���|t[!*��&^�a�xXw�9Z��[;w����Ŝ��� -�ն_ޜ�1���!�s"�8���hI�wd��a@�Bj���JNSL�;| �K'�_S�3��~T!LL�:�؏�P_�W-�ù���?Uj+�ے���Ǭ?�E^e��+αX�z��س��y
T���v7�K:�?G�=-D�1 ��"o*b>���(!��^��b&��������TV50��&����٥f?5	����P�\��YQ����L��u�VʐH��uX�, q�J�q�������k}�l�-���7;��G��<|�E�Nud7��ܭqX]w)���rj�x]��X�T'��(�F?FD�8ӗ�:��݂p��8�$ }���@��.=��kԚy��[���G�بe%G �I���������dJ��8�Kj�,bd�4E������#{u9Y؄�6N 3Q�Mg��͗�ĥiAY��Wˏr�!S����4y�5�Y�q��t��Yh�4笺�������
uڒzfJ�D��r��<wE���>�+P�۵�.��/j(P�������M�$�KE�W��B*�C��� .�[\p@�������߅w�m7�>Q~��Y�V�.0<&|��CW�TW�Zf�W�'��>�B�%�g� �<)w	�T���nt��>�h�� ;K��KQ�*����}�QQb�7��X�p�^��?��1�>�w7վ��/m�5��S��'����ݲ-��X��n8J˝�ƪ���%���{t0�Q���m ����.<,�� l�Z��4n�YD(��F,�A�z~�V�VKp�5Q��̒��F�M,���6��BV���Pŗ;(1�-:�ȞN��:�����5��Ue��r���aX�׃D��s��c�~0�ۂ���b)� �B�:�O4�ރ�j�{n=���֘��[�!���sl��F����玕�)Դ�y�4d�S���]y��9`/ �k|J\�N�L[�n���]�3QH?[��/����>eV��1E@'N?���DxC	��M�J%�U!g���rk�ݿ�������<�������y�ʹ~�y_^d՜n/'s�*A�<��(��@�ڌ�4��� ��� �O@E�_�Z���[�@hꤴ>��mv@p���y�����1$Y��Z�h;���IP��a��<2zϦ+�u���l���n�KI����7��r�u��;����Wzg��izA��@[i��L�>�桲�bVMу��� &��13ty��� g�A3Ji������H�B0���Ru[����'÷�ty����ĽJ�����/y�e&�GH+�#���*�wI��
��V(�μ0u��a��}N9ҟq�*���zMW��9�����pXIS��u�\�`�5bG�lW{��(��:�=�A�C����tvw�|M��cOi86*�IP_G�H��m|��[��ZA�y<����*M�����v�Թ'A��#~JA'[�P���g�2�h��q\�S����.�@��1d �Jl����#j��c֙�����ĭ�H-t�<SDQ���b��u�]�{FX�񡬫�~��B32,�PD�(3F��t�=b�t�E?�7���PKXq���O���J@����r�y�G����>���"�3'�Yj��>��7��B'�?�N�v? ��_�MF� X�\O=��2������2����ώ���&^^|��8�M������g���{���<��8�l��]��4�cy�dSu��ӮM�#�c�P��M7�S�MC.������ [`p�IB�" |et�'�����\r�؝Iv0d���(����s��K�^e��� nZX�l���k��kd���i\"v�>�1�g��q[�,��)����e�k�z.N��c�^*����q�f���$I� K �a�H��['�}��l��鄅� �-l4^��5\Um�NP����8Q�[�|�]�N��sV:yB�;�u|���x(��]�L�-+�W-�f})��Q�_>WEu!�pŭ^�-2��Q;��g=3�)���L��3RP?o?n���W�uHb#�%�de�����qj�h �!��EŸ�c>�m���Lp
8kQ�ss�7aE̬j�������߉��CH�kO��4��^�'u|��Oz�B�:����qY��{a�^�����,/8d���m�sZ�E��u�ϥb�Ll+k�Pop[]B���g{�fN���b*X�kA�5X��_��>h�o��H�p�eeM���A�3~�7qq�/ӷsg�)��s����g�������t�	�>��9�z��˅�E� �)J
�L� 3}��2U��HV���R�
ș��|M���`�7Z�k�uQ�Mf<�����F"%�I���Vw��)#i��4����0�fn����#CW�������HhG.T�Z�l!���]Q�:KQ4��W��no���DB�i�ʶ�v G	�v��U����s:�tS�L�jۜ�+���������ZT:��k�u�$�"=������ȍ��2,��� 5aYWm�CKJ�xQ���!��`%H0DA3f���:��)P���t%Z�άg}a�\�s��t�W�D�������c��W�Ro1�����o�+T�.��u i��.vc�C-�9����(���z�C$��.��FB�����k��a`�Jx�~ԇ�1�y��A|
�D�����ҋ�EK�D��~`9����'f���%if��9p��T�R����;h`�X���.Z	���
$'0Bw�en� \��������$Y�� ^`���	 ��er\����Ux��V̮1pH�K��i��.Jn�I��K�}�פ%b�Ha���
qB�����	���=���e���P���n����A��Go�glv�+�+~_�Q���c,Ș���>�Ǹ�% ݕ&�S5�����Õ�����I������J�k.���.RkR!1�X�H��~�\��KW������F�BB$`�)��{Β�X:�ꄐ[�����MkI��	�@���J��`�ji@���/޳��$$�4qs.��k����Z�7>�<�K+�:���	�<�٫7��������(��Lˠ�j��6b�ī�m6�[V�H�U��<�I��Mg���+45�.��ӡ�<=�wr�Ɣ�d�K�;Q�{f-~Ӌ]��_~ZxC���d?R��m��rD~��Q�� U�U�2�7Pß�K���
o�:�ܲ�w.����
?I��(��:̧"(
�Z�J`6��Ƅ�Po\�����t��9��G�gT�W�
��b;0��u���@��6CQ���̭_����M�V����	���Ã����gy�#�:K�l�г��do �vH	,NM�ZY�������ޓ4^��7P��	\d>�U��ȶ~'UR L�K���r]B=Q�����%6Lkp���٭"����1����B1��> ��E!�j���~l��'���_L�:V'�w�߯�~�3R��oWw���b���dy���OC��M^w}޵��@%ÿ2߮�:�*E���׶]�+�H���h�(�M���P+x� �u�B�;��/���3?���H�#HI���8&�<�n���������˔��t�Ft����
��ftwp7����֓-��Dݴs2h��%L<C�9�C�+h����_�Z�Ǚ�h�Ub�9|�&�+�"Wn�☍\�;��Ѻ����*ɢ��ב�&�}2k��`�\ؓ�p���	d�I��L��}R���C)t9���-�	�g"�F;
zN3i�PL���/3���(u�����GLzc�#�;wm�>���,ga�����[3�/�7ҶGʎp��Hr�+��H�TL�z����,I6�䷙��*N֨@�8�����~�^�za��*��g��y����٫��	��p)�?�
p�^��-9���j��ͼs��D�'��t���T��u���Nv@V?q�[P������uT��3A�^���NUM��DV�����3�|d����}�TM]�V�gtUi��N=O�a_��eg=�܀vN�5p�a9�b�ؽ�x]n0dn��/�I���xk�g9W�^�J�A4��=������˓8�+r�x��6�M�3+�R8��,����P�u\˵�=�j0����*7J2�B�ܿ�&徫B?�_Nb�>�y$=�rǉ�JkabJ^���l���i>|?a��S�H�q;�P� �b̵
Z��f��ʹc�!��@�9��ș�M��R��I�>��@G���hډ<m�W-A����x�\��w�[��؀�E�/v����ʠ�6{p͉������]��h��OL���D�����K<bۃ_w�o� ��ױX�A�|_�hyž޲R��0�9� ��ѓ��®j��3!{��*q_C4`F�Mv�x���_8��d9y�'��s�s��,�4���Y�QCE=K�c4��C;ٕ�J%������`�/0缠5�-k��~lU��;M9�+i�sc:D-_��1K��:��Y����a(���QYY�胉���9O���E9��6ׂ.���kvw����f�Iwf��8�'%�[v����x���!�`�Vpzy�ZS҂���^$���u7�$3'm��@!#��j�~�;��Ꟈ����;�p���#���m|��ע:XJ��Sg{!�
B1�0�$H��� 2�b�U�Q�u�ө��^E\KN@p��R��܇�G�M��N�Ԏ�l����A�c���)���lI�D����"ő/�DM(O��Q�b(��
�U,�=�_��9��1�6�Y�K��g�i	����#{�-�4�Y��:
�'�M,ib*�./��yQ�E3�ֺ��"������ɻ}�����x8�}gl�j�nnHR�E���#u+�����V��f�(�����VoY�ȕjQFg�}� �s�<X�yp#*���9�ڷ�)O�@̇˱���`~��Z{�:�S\�$cEn����(7C۔�i���״?DSNj^v�H)� t�ċ,�H"�ě�h��JeU���U�k�G��ѻ�q��-x�z�%Y���8��:u�mZ�������v���%(�r�
���Q{/:� ���	9Oj��#�Ở�� mk�sMh��������˧�%Id{�xuz:�������u P� @u�|[�%N��Ƞ��h���.��t�=��1�3`}&�9q!�o.Mw��lZHf=皋�G]�S9����������'�CB��d=c�{�eb�cM�c�=���W�T�KT8!HW��@w1Npi�M�si3�ǷҿvF[H�I�%�n�81�Z-lp��ϝo�7$�_6I��t^\�_t��uկ�Յ�WC������_l��1:�zrx��'�$_V2Ɖǻ�h����+���A(�3����e|`����8�)�����ձ�
��q}�e+��KI씍?_@�"��.A�S *^�qT%��`v�H$w�__��Cp4>)Y[�1z��<����v+�1��TwŽ����1`[�k�TT��{�Kz�=1J��ޟ_@�[�:Sɑ��uI�T�Ro����Y�������ނ6�;`�
K������y=�m�]�Xp���B������@UG �ĵZ�&�ڬ*� ���J����6�󛓻nSM�&$&Y%M�[y�}j���<��f���\���D���<8��B�si�F	��|w�=4�$�U|�������8���d<@�_���n2,�J�R��U1�nod	�[���E9��F��`�\�F>���QV�E����P�K��2�ךmt���}�@�N���	(xQ*=P~�u��{?����s �B�um{�����Eo	�b)3e�&Z�7���c�'�QD{����'i���mΟx�����GoJ6��g,ZvҠ%|g�*?5���L��E�fW5�����_�g����?jp�̑���/��\+Tc6ԁ�?#O��@d��h���w�cв~��(���gil����S@�}�@z�R�6�{P�T@�g�tg3V����*��o�$�/_���v��,��~�ʭ�j�eY4�q�����.p�&.��N+�(�i�Z��ɵ뽇��ӱ����w�����Y�|�� �	1ʿ���6c-��"@��(�Y)��1QH��3�ɒ�J��4�@�ˊ<Q�	�#YnS�ލK�בv�.�;��kڋ]�c����F�0G��~~Y%Ij�����|��8fm�����U�U%1Ě��_:�>������e{��)�1��ۈ��l9 ��V��?����Y�����Y������h�� ��g-h�
I_M���Af*���z�^޽sÉ��G	m؀��IM���Z��쓨"XCcttn�Qu_I�r��K�::E!�n�9���>�a�
,>c�����wnlS��j>�t�E��R���X�N��Q c����C�|������8�e���+�jlb�jm�i)G?�a���"����Q�+��hjL���*_�K�$vF�K�L��@ͻ���?�v��e�Tl�n-����������ip�fP���F$�w���Ā\�?Ɉ+e*@3E���K��L�����Ui;���x�V����h��R%v�����VLL�@����y�Z�91���*�؈ن߰�|����9 �a=E�;�nG)� ����
7�
���_~$�7z^r{�b�P��X�=x��)�P�_��b����	�m�Th�ϵe�Ƅ�(���>�y�l�����y�ߢ>#
�n������jsI7����⭶P��X�o7a�NJb����B�ܟ&>/ǰ�����)�U���j�Ij���&��ct¼Iz�k҆|H�@��N���޴jv�o����S����� ��W%wxT)"M�[��h(��C1�9�~��QZk}g�}"�^'+/S��kbn��tSi�jLs~�:)G��ګ�;'{���k���n:��̴���$������sD�32V�d�oU��$�o�l&s�[��1�..��o�{����s_x��n!-p��d��W�ͳ��ފ^a�թ�&U�}��M뎇G*�Y#	Tb��;,�ڿ�ϻ\�>� �� x]h,L����Ag_��]-���5��a���/��n]<�A_�'�t����`L�c��|�K�����5}?>������z��(���������X�r�h�A�en:N�+�����Û�_*qQg��";E��m|i$�S�0J[��7_�ۄ7��.�?�l��%��)˕�PX��)�<���	��S�����I7j9�R����=�m��Xj���N1�^��K�x��3��9o��j�H.���:�d�>�v�lҽ^�-��j�ݹq3k�Ok�~���������0�y����jˆ���ζ�[��N�<�d�J��[����cAA���npk�AD�M	�W�R!���(��R���2���*�t����hK�)�ܮ�B�_�Z����ߴ�;�����C��.�u�rbf��y)	�9�bא%�.{h��n:~�~�Zp�ALg��6{�x=w�K]5���@BN���5%�iÜn��/�dN����>����z��^i2u��0�gb�c��r�c!�UöQ�W�6=W���v�`=�B.�o��ow���q2z��X̴w�{�Z�c5!��y-t����*�\hU\s���AIo2�Kk��_��OTu,�RttP �b��h쵛w�t�������0n-����"��l��s�I�?pW��*^ĳh��k�[���J#L.\��H��E~ގ�aj�1x�'�<�+�}������p�Ixn3}B�����$S~߂�2$��_^ɾ�#�I�E��z]ŗI6&�]�[T�Nb����y	�Iy�"��NPTT����ъ�t~�F?5y���X}�)��;l�JX'#ކ��o�тs=�;�e�D�7��UG��J�)�STUϾ�=��Й��p�Z�tդ���ݯ��R�?�w��FxF�Џ� �}kf��Z�4&���Ղ�}�T�D��2��{�^$�b�M��9�m�	��AI�Z֓ۮ=~�:�0ӱM�1���E�)r����Ia��P��� qsm�
G5�˗ώ��zę�V�*�;t�h�
n`޲���u��χ�SV����.|b�Bk�ϫ �b(N���GY�8���_em��� ��1��%���+�^$��l������'���Fꂲ���A��E���w��]�r��j �b���պ6;���1U���,0@�1)Q��9tl>m���ѳf܎�g�B�&\���������ʶ��� �Mr1�A'�r���Z�����I�]L��%���?�H�s��J���'��	s%���bd�<�$zec����#c9�Q)[L4C2�#k���%D���U�u!�}w�J�o�g�m� v1DW��V�>�2��&	i���s7�����U�̈������:�lY�c阊�=�Џ�8h���l�s!��GG*���o�FOqQ���?2�x�B�4#���]gY��7|��7����K�v3農���B������g�M�Ea��%���i�_����V���8�)�2_��#� ��ƥI��D�1�W��}e᫧:���_��hp�RD��a���@�|�M��S\���m[��@�u	��
�`��)�M_x�W�s^����D�*_:\��8(��y�oC)^}��eͷ�Q��i�޾ZHcDWK�A	@N��-��L�"�N���wr$�>~�������D�."�N?��!��<���
�����:��L��x"o�:��f鄇h)=� ʚ �[��݅�@���R�	Q�>%��#~~�{r�� ;8d��戀��q�w�������
Y� W�}-�}��XZ�QS��5z
d�M!7��'}Z��\� �lT����ga6u>+������������O���s�VcXYPn��s)6.�����ut�o������mV�<{F��z�ա_ �ګ�,�S�qQ����x�5�Pn��K�4]��@�K���.�)k���v�cJ�Y��-}�s���V�Z}N�]����h��b���,���~׾(��v@v��R�sXR��V~�r\��W7[���"wn��ʰ ����?W45����b�� ��ٗ��Z�N�փ��-�/��n~�.=��Jox��3��ɔ��3�wҹ��(% ��++&	(تr�t��]��?���n�����7��)3(v�s�Vc�`�z��qq����f�á��jy���Iw_��;�4�8YX�ה�Z�(?5���C���>{F��?��^AK������Tr��s�9,�����Ɯ�3(�%���37�Ş�4�ݓ[U���#�0�e�w��gcaYC�݌g.�=:��2�(��H����7���p��-���4\!���xk3��M]���/&J�b{zj	{����5��w����י����2{8��]Tp�n�q��ʋB�p[�{���9�����_���|�6RRي��8N]o��\�.�N\MJ�v�H�ON�֫~{�3�?�$�L�:a��>��Kg�;�xx��gKFB�t���?<\!y�>�f�[Վ���y��]�>�
Ƨx�ι��}{�оj[�f
g������S<�{x�)��(k��?cM@��#��%]��7jD�9J�y�@.��k�م�Bm]������F�]�^�T�2.���IBy�7���R�u�q5?n	yU9-cWS��zII��0K{��'���'��n5���*���ollM0Y3�<t����!4
�.����F�oK�G��.<̪���/?D_J�7�X5ʫ��v�>���E��S�'y�ؔ�j<��:����Gl�?f��.�m���}���z�����:�o��,1,M�n%4����.���KL"귶E�v_A\G8i[���r�D�W涺ԅ�GF輸�="z�:��d=���������aGBX����
^ʷ���&?���r�5���8>�_C�i_����?�"�|���z�v��"���Ԛ��3���P�߻JV�{�s|�gU�ľ�[���p!#�c�N�z�TH�v��1���pm9H�v�B����AJ��#�w�,YzD�r��K����Z����Jb'ٽa���-r_�o�~<��`SP»���-�p����x'>�ɲ�E�E33潊��rΨ(�ƭ'3��A��lW��C���X��ٵiji�����H�[�Ė��Jaۺ�?�>WX앞�w�l��Z��D�T�<-�_�*V!�i	Jmv��m���j��t�u���C�_nT���'Y��mM�ꉂ��g����>-����Zפ�x���_�,�O��H��|�o{/�b����L[���_��<"�l��'?�˾�j�\M,�IQ�s��s��~�Ob��U<�M2���A4~�G�Pa���#W��F�ޅ���w�%�����%E�ƅ��������x���p���Sȍ"������m��C��x��4g�l������ϛՈ��t�oWGc��#�q:�D|v7����#�"�voI�Ռ3�;�b��lz�N�\ˇ�/�O{���ń5̣̜�����mf|�!�Ac��=jtB��>��j��h��־܆s���y���KT�R��q��MfW;�M�m!�T0�Z43:�V^�^aQ=ȦT����8we�O�<�e\<��(����}��5����|����u�gK�%��E�=(R�Ԛ���bW9�}-���6��VZ��Yb��g�k�с��G^�ֱo9]g��S<��H��~��j����h�3)ɫ����@(TM�	��Z Xa��"a�_B�����@|Sb�.Ņ)�6~m���w(.�m�X1uxL����A���џĐ2�G�FZW��?�O|�7	�F��?�U�&]>�sv�m+H���I8X�w���?�FtGe|�}�b�/�����F��_<�3lZ��*�/�E����r��<�Ɛ���K����у�=���D��6��9��o��v����j�Y��cU*�)�oz����ډR-yE�f+��3�zi(��X��_��3��ok�&?��lY3�=�Nd6�t�L�4��޽M��E�I�?��Αз�J����ixX��{�����z��$�6R���[�4������S T���Ӵ���KU�%��Ψ�W�M�Tx	,�� ��d�e~}i�8M��(�O�P���hG�	�1�d������{�$���F���u������7�)�1�ѓ12�E�=j�l��vzq���>*�u=�?�%Qf�OL�lם�c�<@���?�]�����<���l�RG^H���v4��t��3-vj���tq�n~dM�xh��ɮ.���pj1���Vt+c��L�4G:���sc�k�+{����j����XQ����8�-Gl���m$��8��l���v|eʝ�����͕���:��#�f]@��A�v�+	�}$(E}S�=-9A���66���۞�7;�20�W^%�	m��5g����t�������?��l�o�(IGw��I����P��gr�9d�o`2�'�7r�c��>��-]�P·���^c_`_PA(=��]���c��:$��͛6"�YE$|�ͼ���!gb��׹$JX�IND��1�u�!�?��r=���7���5�+q�q�s��[{۰��g:��{�A87����Iv;n8u�՛��uϓ�_�M���>(j��h���GzsPo�fl���A�Z	
��ƩT����������ݽ����o��z��?���P	݄�N�R���q�pJ�ZH5�r�Ƙ:��D19��\Ɲq)Br�}3B��m�����9��k������}�?>�����y��콟�_{?ϳ�VLٝ����*.P�;0ݏ�:.����FO'��H��Da���`F֩���͟�u�\��I�J���,ª����&��o�t�4���d��U:�����:�[W��7�ݲ'�����ډƇ��i;�;>&5e�C�'�'��zm
���F�k,�Xg&H{�\�C�~}����'�Y�/�
5�I:���c�'�Iϩ]nM:�i���h�$��@pAn]D;_˳!'�O�l)o�LUG˓��RU���ߚ���"�Sfg��y_@UJ���h��NgE��/�������'��E��gwr�����x\���)z�5P�'ڢ���y3V04���.����dX�]�h�[>k�컵G�p_����Lf��yJt���Zϯ?�4F8@__�z�?�vK/�`���^�8��y�A�/��o[M�%�(��Z5sp�����8I��_�2&C�����2��G�h
ޅ�s�g��]���ۍ��>���Ά��ϕ�� ��]5E��� b���&��������a�|�̳�����CPt�E�J���8g�޲��:���d��u¥�@ae_�Ul�ǯ$[��?�����\����}��t���F�ڌ��O���ࣇi2�"NǨ���UA�	�Llqcf�v���#��NЪ"���+�n�<%ҫ�׹Y��g����y'�e5�>��^uv��YoO�h�&���9���{�c�Ǚ&���\�oY7.�\p7��[���)���m�������7��Q�98��V�ŗh77�^�3��um�����g������Y�^p*�mK
���	@`�~�}�EX��~��>O�+}�Y���IbA
D��2s2�������o2O�y>K�P�`��B��yv��EJ����[ ����%C.�����h�^����0Z!k�CL��I�ͤ��F=	f����_���cw�4S�\���'���Tz�'��'�0�՚G�ӿU7�o~� �FS��^t���X)7c�(� ��U���k��,�[�Ӥ�+= ���`�F�דB+���D��t�v�?���|@�ƓPG|2���Փ~��SƊ)&���{[7�"�@˴8�(�c�d���O怈�g�����q@�M��O�Y)>j�h��H~T�>ɲ艕���"a+%p>�7�T�fr���QRt<�Cz��z��{��w��o���~s�K���ۊR@����wΒ�4�[�����S5�˳��5b��i���/�O2��^|������Tx~T��Fd���_��-W8���z�u]�Q���|K����I��hY�
ώ_n5�~O�T8[8�P��~z%�T�	n*����� B��B,����`�f[[2く$ō�hy�������c�j��)9�����09� �š6���p1��,�1��ͼ�m�/��^�nlf8h}�������V��t��&n��~�|ŉ(�ɪS��Hg���xxc��s!uN���=�ƎE�v|�}�9����%o��?L����ݦ���_�s���!�{O;���..������ڜ͵��7�z�:P����9��=��=-��'� �jՃڳ��9Okt���aߌ���o�l���VJ��������v&q�*�|1�χ�o����~Cm��L���"F���JF@N�e�1ӑI>x�ox��s��������hw���{i������K~_7�7���k�δ����&���|!S�Rq���\�|��,а���*l���ϵ늏	�K$���*>�9F�5��>�0_�G2�/���G\��ʳ�>���Zڕ�X����L�Gd���H������I��N���;���*ߖvfpW|��4s��������܇٥>�أܸ�������<瞄�ŮN���m l7�6�������J=�_qk���"���a�ƧCS��L��~���)���V��ǡ�M)K7���uk�~�>��큨����^����qt'}xTK��usa\H�Ю��J}Ŷ2!N���`C�R��(d���hE�?��՟!a��q�#A��[�K"��7��;��� G��UT20$t�wxR��}�r�r�s��m2�t���i��0k=�px�ϟ{�)v뙗/����s�(���K�C������1q���e5_��O��}n'�x�o�X�����<�t=LD"X(����Z���K�O�½�i[��g�>��$_�&�>��l�a��%���. r,�b��2����k������l���}�����ot�vvޣOyf�w6l��a���Yh��"�M>M9�_�P[8�Ԧ�DȬ`<�=R��a���x�+ ,�7R5���fT}���#�xy�;���cJ6G�M� �D��u��'&�/�,�����QR�L��'DP��n��D�ٚ���|�y[k xW�l�����X+!m���(��i ���ތq�M��hG���zN2�Iwj6��x����Ĉ�?z٩�g��˅��?-�SދAH�5�l� B�3�1�����3�k�1NF�Ue�.H��L	ءj�\�X- �ۏn�p�yߵ��n;��#��������������4�8����U��YӳG�d�,'����A\���Gt-��x[|��R��H�����﵏0����/�v5���9���P�E9�����P�>��X����@b��^}�c��IC�ӈ�$����������+���<�F΃�+[72��l�0��
\�a+)�ux��e�m1��ƺ�u�h�[��L�Y�XM��������ӗ��3��k�Z0f���C@!`�S*�A+����Z7�g��,�3'�ioUS*��6/.����؋�>	��}��f�K[I��?�"�ɍ��a<~��ļ疵`_1 ؆�U�4�n��)E�iuA3��$=�+6œ_�B9�#C[�8�2Iغ�wC��ĹsN������nss�P��=�X�@�A`X���S�i��'g��{_�Bj�UB'w�ί���]� @4?�zB������/�R}\�A}5Ҙj��o�X����l��%7��{BwpL��m��|�u��r�6&�b����`�UL�Y��_����,PnL],���L�$4��$�o�W=�9e�_,-�?PԀļ���WuR>�V�� AD�Y�nA���P�X��ԟt)��Z���i�4�DJ����b�ߐi��^}b�Wǅi�a�����҄I�M�"��>����R��<�(w;����	w>;��5�w����eeV��D�����{�d��e+T,h�$�	�:{#n�6IKK�)����B4��5����5tjQ�@>oz��}6�$�RxM,w#�5(?ϟ�F,�r�Mq%-\B���>��s�wFNB��40�չ'這�Q`�L�� ��љL��C�V�
dV��BZu^�Y�u}�O�KY�WCrZӆ�o�]a�''�o�;�U��Wjv�:W;t�g�Vl��FEn����ԴND�Ű�<�[��S�g�kX�X�)�n�ԛ"�+k�^��9O�..+P�f~���s)��ؓF'C�`��}��(��6*%�������u�t�O4��t������ɚZ�JZ�[�7��U<�E��Ĺ%!���f���G��PEfN+�PI1��� ��4:BҀ#l��(��$�cf���5a^�!-�B3�c�|���{��ú�F��ʗ3+G
���6C�!�tZO���#��+���Å�BZ�<��5:�Ҭ�75�|��� 7��C,�!ۤ ��҂'G�#���<*��d#���A��.���%��#R�
<h�l�ş/�ѸXo��}!��xmh山�~?f������j	�K���T���L*N�Y�%��0�k�'\�|2+���h��3���ڢ)��Y���O�G���˚�WlZO�8>_��j��~Ya�ƶ��_zA��yV�;�����[s���;��{����V�j��g=)��Q3�FJ`%a��T�G�kV���Ԁj�H���� �5/��DljW�}���(���%2,l�	jω�Z2U�iB{���j�$T���wz�F�a�#^j�Z\�8P�w+��Щ��Ǭ�=�����}��mJx�{��O$7��ܨ9�bpPF���X����f��{��O=z���l t�n�X�MǨ���кɯW�9.t9_���"��B��ǫ!��n���9n@GT\1tm�����i7���V�D�nB��Ʌ4��G���H��\�
-�3׌<�-�.�DӪr�����SI�������)��^+�����,4�{��f�~@\;6г�"'_l�v�#�
ǫ��`��DO�z���;"����SRܢ�
�rm�w+�_E}$��yl�~����ۀ�����tsV'�w!#17N��j*L��oK���"|q-��{��>�>KԶ[Lc�����S�T�]��R������˚ׯ�`F���dq�����JB�>�D�)B��:��4����!�c$DǓa�(� �ɳ/W$V-w|ծ���YRL���]�矾Q:R���bU�7%�L�+�WO�
��Q(o�R�Q99�~��q�Ҹg7�CZA��Po���)��v}y���Z�rO�)"H���+T7��V�Mm�����˰(�>�+�`R��o}"&�[pK=�Ӆ�^i���L�d��0Aǟfe�3w�:K=�-�d��I�[��e��E6!!��sH�kT�%��� �5fz@�P�*Z�8�<V"�A��Ʌ�6E��y��\��KlZ��$�:>��R��a�nn������Zz���7��i��X?ہ�� ��d�!��`gٜ��ѭ�Z3����(��>������q-�A�H����%r\ͫ`|�^-Ά�{�&T�_h�9:FS�Ѭ2�(�G�C�mW�\��c�����f�a�CT�%���U̬[,������Bl��R/SV��]`[� im��]�>s�Y�%�]S0��R�u�kOKG^���(�Y3U^؊��M	@Ϊz��"��~�ȧ߹{W�ۘ���Lor��!)�=��c�F��ӧ��iXx��͔���a���ѐ�N�}c+��b/� G���� ����`{V��2�|U �=�Ɨ#�6Y��u�2��~�)`���{���/�߁~w�7�r^��4V�E=��_�%>p�YX���?�c��� ��>0������u��}��3E�w���afE�z���kR��_��?���C(��l{���S_������mւ��unF˧�O���u%��v� �.`F��� DM���^�%���鋺CĕJt�h��{�lQ�SW>��Ea>*)�����c�==��}2�����|���as���3�tm���aBF-ͫ�xh�F3��b���^���ga�HXt�~�p�6}��9_�#�g��ܵ*%R�˘B��R����ܓ�(�b�"�Hd$�-����@�:��u�jJ\�����|�F2X1g�3W�}�2�HV�;|��9B�p�c�I�TjO��f��Q�7A.����K��~]U�=C(�z�M�R���y��y*�	���\Yq�l
X64�3��!���O��q����琚�W��g|j=Vuz�%�؇��,�����҃�3����L��]�G��3���O��T
��e�y�ȴ��.,ww�u	�<�y��	v3��ɯ�:Oɻ�T��t�dV唴����罋��u�dn��,a�i��ʩ�Bx��e[�b���)�;�RU��*_�GP���Щ�wa����>�Y[l��`LF�ɂ���Cuم���l��k]�S����0��#ֿ���3����)�����T��1cp��Bi�sv�r�?:��Y��������:���!2�j�Z�u���@��/�I�i� �«�4]��f؜�F����Z���U�u���ԃ��o��'��3�<n8�X}l6Џ'�����_t�r����ċ�OXz��_��M�^�׏�su�{�7v+�G��(bkk{Ğ�|���%�7l�~�=0���{Vvʜ��� �����J��y��^?����zd��0&�o�`o�s��TϞ�U�����b@��N��Tw��n�MJr_��.����M����u�<���f|��v <
j�*v�S�޿C�K�4�q\�:�8���Tk�K��{��}.��Z�)B��wq�F0��Yr|�c�]����
X3���gW�m������<(�[��E�h"Ǒ�{�^Y�x��V�W����}��<6�F�C�x�"{�i�	Nj���.�B��J��4�����҃�е`
�2�!��xSWd��^�e�6�J��>�,B�^���8�'M6F'f�5%%� ��{���[�o��#+��؇��rət��,���ڑ��+�'fĖ��6�N��q6@�����"EIOz.��,ao�b@��q��{�4R�~�?5��4�,f52[i�+	���z������Dƫ���\�}X�P|��EAa�OH{�P[/�%�	y�$ ����&�!E.̍^�ڡ뢑|!j�VN��YF�U��}��s���\\5H����Im��I7�SS��>����Y��&H4n��-���n��Z`2}����%��κ���vɁ
���1۩X��v>M�rt�H�w���n�7	C0W�h����X�ʑ�{����t��3��?�������"���s-(B�w^�<��vt�S%<4�0]}h��D���M�X����|ĵ�&�T��h���_�%k�������l��I��0����=i.���\��s���`���%ȷ�����$`Z6�TU��"�X�F�V�m���i�|�F�A/\N�&
:�`��TJ�}� �}T��Cb>ח"T���&ȌY�ݳ�z��c��^���D���]�ri�ң#& ���Gh����se��7lN��Z����vJ��s�Ņ� ��Qo�x� ����e64t��S� )z����Vn@z0��M�,D$M��{�������ޥ��1���X(v�ц���#���^�۾�%Rb)a�:��WV%��mY�����-)4JA%� 0��A5y�7����\V�8�)>u��(^����v��W���"���@jV<eb�>ء:�Hzj���`��j7�F���f���1�E-�W���U�E�1ʾ6���Y�>[�}�E}�8i)�S
3��^fq2EØ�`�8��pA@�n&���}|դnw+e�V��J�>�}�������Y!1-9�s�& ��Z�������q҂.���+�\|߉��41���>��؇}7y�,�/D��-�D�5�f�Dqx���9��Q�� �&FNZ�����`�u߿eG(�X�r���a(��l<�����F)�V��G�|���ZJF�%v�-܁��қ0Nf��E�C�U7����k�)���.�	���g��z���+;$�k);ʁ��^��!�S���1jb9)��)�>bJj��
�grD�����Oos�Xo��G��i�:��W�����6z�73�jx3����>�?�e-A�C7B ���b�7���J���i��\$J`,����R��k; ���Y���S ��s�K�E*hҳ�@�\?��V/|�uQ>�x���{#<�8"�1[}U�E�`$N��E�� �g�@�{1_��z�/�]�� ��"��i/뇇+9����,�}�*����R��M��e�a��c��5��Z�
���'❵�Uv��n�ӕ�A�¨(��m;�Y�0�_Kz�ѓ�F[Q��:Q��#(gzx|��!{Q+���=���yxo/0w//1�▎Z?4z�������'���dqi!��D*���mr�:�ܴ�wD���&&���k��WoK���r����63�E��,R��rn���c��͝	�=dN3#!&�n�@W����b�����>�+��S<�,;�]���^�]�Hm ��r#�	[C���3ZJ�	>�}�������$_o��jh��[P���I2�
�4����_f�ZG�o-��g��Z"!��^+����c(���^�R��ǣ���9i���]i��[1~���'����]�߆�g���7�	������}�l�qm�'8U4�Gk�~]��'YA����5��e�.ktz�\��!$�U��o�Ё���'��81��]���g�ֈ��J�^���C���$EkT#�k ���a�������l�-���T��Q@�Ĩf8�em'�u��~���W�S��)�; o���S�̛�����1$|]�����`����f��=�y>T"v����4%�	��_�2o�e��bz���8(��I��v�ˍ�}�/��W���G\ ��D�yR��L�����m}��Yk������l`qT�_�(�����4g�'�c5��$j,��(:�e��CN���ڏ9W4S��e�?&(=|>;�d����N�	��%��oQ��){\,�V��8���o�:˂��8����]�q�T~n�|W�"�D��M1�l�!s�Ă��'&�ɛ����E�r��9�F�e����:^]i]�a$��@��;�yM���dh@� `�m�x]*�X���:�q����o��K��U�R
j��S*���4���5����]��oUi��;�»��	����x@�Z��y`L;��4��t�A%qT��b�����D�j�t�"�s�L�!��1}4a����`6����ں�n��\D��j��I}��qك�[�u'ʍyC���S �^!`�^��v�_�Ms��N�%Rx�U3��}���{%�(�d^�ӏ��ij��7�RS�X[�b��U���m�P_
���������*�[����*\T�<X�3 �I�*���9uX;`y+ሄz=��I���;�{N��H����|ח����|��u�d��G �t�'��T;$E�b��D=���8�	��+Y'�&�e�� ��9qq�e���	f	���`���gR�s][lr�����f/��g �F�z�� ��a��K���0�P'��~샧�Kn�X��w�̙i��Y��S��>|����v h����*� ئ'tPE�?�wݙD�������WM��-"�[��x�s�p��]�������ѯz�}Q��;���Q��	��=�ܓ��B�k<����rg�fҽoT^�����o�^� �l\���2�U��i{�g��R��.�=9F����#�e�R�Mˑ�T����/1���8����y��3�E!�ߴ�Ij���uj��h'5�%�GCh��}<��HT�y�� "6��v;`�Mno��L�N�8�W�#3f��<"����$>���W��*36�g`���i=���s������
��;�}��p�d~���>���/�X�ґ�#�Y�9෥��H��W�۷\7zntspEK�D�-�)��y�F�v ����j��Sƴ�X�76�HW�e�������\�G����v���7��7m�����n#_�\ch��D� �(6ࡏD�e=4����	��3w܆4��3~>yl���F�3�9���&?ieluh]g}���`F5�[ۛ��(��ۀ�����f#<N;Ǡ�d�*@�a��Շc�Ѳ�_�� �B�;��%�~uVr���?w����"!O�u����u�>ƋH���;̶d��q���s��6��7����2F7G����>����G���3��TQ}V��1H{EP0�����n�[b��(�::���v�F�@~�){�X8��g�A������04V�5q�:��ow�\�Mֻ]��I)"��:ڤ`��C�D��8�ʛҜ�R�����5ЈQH̰�޼3��K�Kqr;�^�0�0S������k��<�q��R�K���s'-�NA�S����5�þ�7�3��K��ݤ�X�t��Ge_�J4P���U}���jFʣ��G�ň}��:��v�%[�Ja#0W�"^�*����7�a]Κ�Κ#�\�F%/?��MΥ�����=A���:o	��<:-�����ژ���Gci2��`\�|ձ�'�{�D���Gy_b=[�d.����VD����B�А4����������1P��a�r�S�a�`[�Pp#!�Գx�Y�~�$K��3����-��̓�Ԩ��H�� }��Dzwb��m>�O�/��X�q�X���A�/�t$�f����ai��jC
�|�����2���(����u���;���v,��JY{m��.��|b���4W�z����}PaS|����A{9���Hj�9S=��d���xܰ˸�ĘZ-%�A�L�~�86���ߗ Z:�au�5�w����m�tC<݂���v�p5�v�dp�*��X��C�1�TQ��v����'�.����������o����E!���Щ�N��3��D<ץz#7�����6�Br��yi m�w�MM)q�5�y�H1��l�����Lp�����T�A���:��+�eG51H�?'��Uu6_���8�/��X��9�t�`�Snա��	�XR᪏4m������� �=!��F�*�Z�6�<��Q��������,r]���r��52��߄�J8�G���=�$MDѹ^8�������� �:�aX�My|����z���
ER�]���W
��p?���o|_�����k��:*+h�OJ2움���*�@�m�{�~��+�Ƭ��D��PT˸/٘s����\6���^N�2%)�.�q�XRv��Q&:���?�Q��DZኋ����}���_E�|V�^����?��E��[ p)�y��;��d�*MØ�1�n�؞�����v�ϙ��4��qJ�ӻT�sp��|4��J��	���V�fn�H\.҃��jg��_\|�$��?�rں�0�m?/a����}��^��h�ƿ(��t���k�志� �I��']�J4H���;�����jo��ŗ��'�-�]7MU�Xz#LD��]����mZ}�1�!S�J/¾�`��{� �[m�?th\��� �ɣz��=���}3�]�_z?6GR���f�'l�U���������k��7����Пa�
���[�A�V���ǉS���#�A��n <_�0n:JT���q�I4�+�Xd+��i�.�xa��2H�BQޓ�X#}a],�����]��=#d�uo-kݸ��vK<��$�j�oi����xs�6�=MbQ4l0"��k??��x{��8)�H��C��W_E�n��%���{!��/o��I�w�{��p!���&>53��>фk1G���,��i'��7�6\4T|�z@���\Mx��&F�'N�w��ðBb˗���h+Iɽ�Kwţ�<�C��׋ݒ��eA L�^zw�T\�܆�ҟ�|���˫>^�P��\{z���8d&.��nMP��������(d�����	���!O�\� HEU �w�/�ﲯ�1c��P�}͞���CQ`���!D����1=���\{㑴e�������p�hq&I��0�}�� �5��J�eL����k�Y�2a� מ��bΨ	ݪ�_)?j5�;c��L�]̪�`o�I_�m`H��b���	����1*r*��j�[ťh��V",S:ڶ
N��*�݌k��V�HDJ%���胦���H�sg}җ�˔)�:/�}�ʦ
K�ݓ����e�U,�Q�H����Ef���x�gJ� 'e٩��<���jЃ]�������`įu�o����n�����3E{D�*S4o�������Z�٣	��r��}��	�Aفm�P�\�y������YK�,�x�]%* `�tg���t�����X�¨�5��(}2O�^Sai�Z �dيJ"��8���"{QZP����0���2�R˜?G����e#Y�8U�m�:��s��_}~�Ud�'54�^ ٮ�L����S�&N��2��\�����ŷ��c�.���f^cƷ��)�Hs��M���$�z�h�y��M7C�E��qR�<
�q#IƝ1={�`s��7�],p%3���4��v{{�,�r�'��M�'�	'.���F�+H�к6�a؊�pA��Y�ڵ�3U���>�o���1M�w�G�{��ٶ��Z����:���W�e��~�J4j�'�Flέ*ܕ��U�\vE��*���U��n��g���S���½��ى'$q��|xF�ڹ�:�J��f�VuEF���w/�Wĵ��h{�J��WK�4��Mpu8����g%&��$��vfA��M�1վ��	��O��_�`��&&G�F�*FH�$	��|����H�x���>l��ths�1�E�W��4r.�S�E�CH4�@ܩ�GG__ �
��"!�ta���Ǵg�ܶ8�D���˗�V�L�卋���$��,�-:��0>��0$W����eCܫ�io�z�9d|�m����hCJ���B��L���	�P,�_��.Bs���t��kĩ{T��8#*������۰�ZZ�6@���l<�WѠ���Ky����p��}�8�X����~E����"ި�<�y�V�_r)a��zU���bo��4Wb���`CS�=���3=t�KZ��;����n%����W{�n�C���ӹ�2�UA�կw��R�N.i`�������֣Ao˽�߷}��Jl�Ԑ��Xh�p�7�ё�lK$u$Xu-���ϖ�@�>�):C����B�m�C#��,��ՆJ���x�i�HE矛���� G�9G	�&1���#���ݼ��Ǎk,bP�[1_���C_A22�n����ry�e_i�!�e�}N�d��
4G`}�"}���J��������6��mR�Y�m���/�Z���àU�h�rgGY�* �j;m���їL����Yg��*ۡ��-&W��D�\��!N�}�U��s�� 7�h��o����@f�ZC�6\�.�w�h�o����&�4§�W��v��##��
Y�c0t���Z �Ԕ�i%E��PgE@�m�ކ������s�O�⢉��u����O�v�؜k��<���j��:ۉ!���]�����!�F�Zs�L�gW����d��q�BJ���Z>�<-�!����0L��0���b�۪�Z/B�%��|�O������>`�� \�����76�喫'm����������K��y�g�@wF���R�)t�^�5�S�TO	U ���a��Y�m7��R^;-�Ь���T	�Q����zH�Dq��B�]Hc^�"l��f�O�^�Z)�cya�G{¸��B��u�Ĵ���?1�ϑ^	���,2V�C���n� ��.���Mz��sj��=�8���P9sꋾZ���}=�U�q7���%���O�c� �c0�=R{ч����m6t`5���>����:�����u�P���I�2��*�����N�b=����H��v���~rɋpibǗe�v�i�r��Z���b���0�� �yqV�݁S�d�r,d��1m���҄{9ֵ�DZ(���R2�,|\��ڒsc�=�V���dO�w���#dStj���h�&v�_�}Rk� �]W*����ۣ��/�rO�)�E��_�t��P�7����a��,�ݟ%����&Bn�~N7{6?��i9i��;�x�o�ϛy��)���9T���	�[9ۘ�n�Io �@��� v�hZu�_@ j�(�3�j�4O��u���ȥ-7'	���+�}���!���V)��5O�b�{��uV"��~d�3N ���r�z��ί�Q��#����В������X�nx��(e�s�7�%�?��P�IW&�6��;��қ_έ�E:3�=�8�꤬���2�/4_Y���ߧ�����׫D ��}ޠ�A�h+;��t�Ѳ�E�X@�m���	9�1nP�?�L
V=Z�����X����Y����W�u��x�x@Ơj�kft�j�	~y4���z�ex��.]t����(w���&��+Jl�����M�O��]R��q��R�ĭ��7�<���6pV%��������G^5Wf�M��)�ϬT��Y��2C�Da5Z�J@�dP=�z�33���z���2Kmt�m��k�s�B6=?b�����V�Ikc��&%V���3�H���+]��Z����%3���:%H�z�ǘ�{�A�G� Ys�#l#�2^�#ߧA棲���C[�N��j���� �NʃQ�
�����iO'`����T��{�����k�=�g�f��sfx-m*$�`�tn"��/Y��ZWE9�事�PGH�H�x���YP����w�n`Bt����L=�m�F���^��~�HHo'!%��49��($��P:sT�������L�d�͇�͑�݀���PG�̱����+���V����=9��t���+��`R_�R��zs���� �'0�`A)V�[�5��ZTd�Fi���������� ������X��^��|��e�OԱ4�������9tBy��f_j���T��{5��)yma���x���������s}��Y���f��Cp�9/ׅO�U$�������01ƹ�w]E/'Ӆ���ţ�H��U;)�4���b`�
�i���f��|�X�g��PX0X� ���JCم�tb��g�c�-̺g��n%ƌѬ���O���.��t��I����)!���>�k�{��7�h�0�ހjD^�C\��qx8�tA|�5��	���H����#1��F��iɍ_��YQ���A�L�^��`��B_G-e~����5���_�Q'��J(D�m���<��Yߕ̨pk�%����e���uoH��?���`�2���fφFN0�'�Nm:�8.@FP޾�H�wG�I�H��Lꋏ���}�y~�U]3R<66P���J��_���,�f8��J$��H��O��*�K��sL
��u�=���g�5�	���wc?�\s��h�K��4Eь3�"M9��������0�l�{��w�_ T^�t��LM�v<9���')�8C� �I����'e�f���'�|7����/'�WS� 5�P���YA������JU:�^�P:{�T1,�A͝ȒМ�(��$:�o��}��b�O�P|����`�I�<�b$��˕��qEE
��aM��77ш;�H4���)iR��p���S�qf��0��Y��+��W�F�%9�(C�ṫ_�t��ѿ����	��ōή��c�-QW��LR�x�c�ל��f�ƕV���9,V*p�'-��n2��݆�B]�	z	+�f�+�ޣ����b}*�	�=W��Z�=VSR։F��h�U�q��
���K�ߪ^��*(�?��E��{��ĵ9yj�K##"+�.J ~%)ZX(9��:"L��A4�$z6#C~_wwNBy`NK3G[��:p����Az�ii. ���V�͖2�-ZL�7-�R����Ou��}h��sYX�}���s�ˍM�����*�>t���Q'UP�a�\`m\�s��te�PJB@Bش$e�.'�i��t^d��c����\���!�D]w�VL��ޜ,�|���ׄ邗��{�O�h^6�+A
{y���\}]h86��U�h}hD�B�4b}�t`��8�MO�ֶU�������i����t)��R�%��Ғr�{K<K��྄��̦��7����jD�b=V3�9����l�p�2��vF�ЕV�k9wlT�*j���GA��p�ݭ�s
{���p�bX�D`�0K��Lu.�NV��C;�G�����Y�0.�ngM�'�s`|�T��f�V���kgBg�ӛ[�Qw߻�;nP,S:"4�p�6՟������	��<�t��> l���X��zx���ˏ?�˫��߬�$8D&|T��U]h+�R���l��]�>��x�5v~��O{s��|v*�Pws�j@�y,���*s��G�M|���snO�7Xh��ʾ����{�J������y�����[ <B����L���* �J�`.�Ǌ_J�.�����,�>��d��@#��G����Re����0p�@�1$$���h�^����a�U�.'�n�9T>�G�A�GSwi¡q�.���I��$/�? � ��i�����P�x>�S�$�z;�h�x+:_u	���x��������tb
�_�v�G�q�"�8k4P)	����HxUF�m����wO�X1Qb��Y������v���GS�M���ͼߧ���mJG�����i}-�"+|#9�����
�;+`Vn�~�>Z���l�WOn�.?.���u2�������Vɺ�J0�H�N�)"�����;Ds���f��9`�7N?�ЅZZ'�����n��[o� a?h�0�*������h�ޱ�B`�
ޗ�=��t�I���4�M�������k�ۉ-V�=�Dm�+qA��	��W��O�n���0p��K�/��4�������]��� �}_�@��*���1��5l*����Ƃ�&ٯ�f��.����*k_p�@,��ۉ����P�+�g]+,S��V��Q�>�Iqد @k��F�/E�'v�%�u�N�գ����9�c��O��cLf}��������ߞ��9�]���/�Ɠ�{�n�������~Y*������#ɢ�*`�D�㼔�����0��d-�M��Z7;�����ߕ�޼� �?��c��tn�#�>s����l�ވ����엞��Y�7Ȭ}5Ij���_j������D��ٔY����2�0c�޿�N��������|��]�ީX�T��RV-f�������o���#�ϰ�-þ��3�F�G�$�e5�T���?6�������6W\l*���*�C����/����|#��ߏ).{���>�տ췶�~��ҩ��N�ߊ8���3�5�g�e�8l���5a����N��i�Sn�=�ߗ��������+�~�0����=��3���ϰ�m�.����m�����ޙkn��G�r��~S�s�7R@e�^��(��ݭ�W�V��h۟��}��T3��g�E�珋)�8���s�"�mr�]Vd�|3ӇpBrs�)��q(���3o�w͗$9�M��F5=Mj���UG��8��������ًp����rox6��Z��a1�>I�r�I��,�Ň�����F����w�W-W���&��pO�zj���j�Ղ�$P��N�#�Adǒ8���AA��/� fST����g����^���<�ͭ��y����xT[5�S�TE�SϩVklQZsK͢���O����Yh�h�1A�UR51��HB�)��i{�{}}�}�+�p���k��Z���p�=�5�@�ը� u]Ǆ�LW&���t�8Г:�[K�M����$��mi:��ޅ]<��%6{�_��lȵÅ�f]r�	�F�qY	��'p� �.ߏ�~��}��ZC�;�ډ�ۉ�3>2A�n�����]#am���ƹ�O�z�|�.+�P�Jb.ީ��rH���Ύ���:7��Z9���o�o��_j{����	�_4B�gu����Φ>L	l^|��d�}��������>��@'�����p��yz�%'.���[��]���_�k�Y7�d�p��|s�I�XfR��L߷n�"��YꥶE�Ie7��n~9���5v|�e���:�Ӊ��9�7�K�/��O��<���/���#.k!��뻯h|��O�Pp�ܔ,p��喽,ʓ������� }U��s�^8�)����lqs~d��T�?�w~kOK�|�Y��T?�5-��d߼��������ѿ�\�%��
��.����(I!�g�T�W��^�h�e���������VZ�S�K�A�d���]��)X8^�2�,p��xWAA@�&�I*� �VzA5_�ۣϾ��"l�L6��T�oW^}Ex{l\;dg 6m�#�nO�s{��eZ~_�z}sƓ�A3�99��C��HF�S�u\��|�]r���﴿�h�$I����g�wc�m_�°f��-�eT����vR��>�_��ƈKm�oH�CS
�b�vssË}��3T��<�j�����[�@�Z|3�T\_�������f�� ���=9��Q�	�/�WB�D���́[)f�\�q�]�Y ��^�}�S�����)�Ņ�6(|���%��ϡ�߈+^ߦ�[������/��������%�V����@�ا�jt��>yr�V��$Ss�RUk����m��G3�Tm�ۇ�U�J�>����%DN"d͢?���KY��֟�s�FS�'59JSDX�<��C=�C����ӂYYZ+��И��	u�����E�A�o1�d��'="�������w����?Z������T���E��*�փ���K�Pw(��5'��]D�sq��k���"��]}iq�d��Q��k"��5��lB$G'��k��؞��F���fA���ڵ���OgT�?yr�l�=Ҧ����$NR"[��@ou����}����z3�z5�,�U���}���\�n����Jq��I@�tW��Ї��B���?�+Gy;z�7�+�Ԭ{m��cj��@wm���@������`���FbRO��Lμ=x#2+*�㇟���Y��&��Oٵ��͠~Zq�jt��уS��f��=~IS��A�/�=�}�H���hE����M�(�C�'������ٷL�� iZ�F!��[[��jo��e����j��Y飊dղ	W.)�?�������_�dYA�`�Sc�Uo(��m��qO�,�ig��3z�z��/V��m��TZZ�4?���9�U���$mhB\%wHD��%b��{<8�m�\բ'�w�tlpr)�3�����<�01q����~I�"���������%�v�τ��1Et���}W˺��?!s�����07�di3O��_��W���`j�f"ȃ���	�
�26�x���ʒ:z�;���4|�N}Ig"�=7��Y{^���+����_Ԉ�KU��9�X����.8����T�t��r�c���R%,�P)���@�5�Ώ
���m
��TM�uɹvpZ]�� ��⭍{Y�$��waV0`)	���ƒ�:X�Z�sC��s�hO��fF���u^}�=�6���R�I���¿ݤ��ǍU�������b�=9t�J=�v8HQ�B���O
��q�E���=�[ex���>�Ao��t1|��J�5G'l���]?���I���$u�����������������v�>x�@[���&[܂ֿ�9��mM����v�����9i�u�u薆�E=����~)���3�O3�!�hǱ{��䛥v6��z������%�%�����	�Ծ�t��n��E��>U���`W�p'�IuX�$a,U��)t�Č��Dg�����w�����=�P!K�U��$�M���F�Dy������>��=�S�I��k�c�S���p  ��#�oe��0a�	#L�������@�ܸ��hJ��/GН���c9 ��5@ôxH�<���8 �H����C�K�x���ֱK=]��'5+?^��џ���w����������DS��ScfD$�|��������;m�^n�aǋ�K4�?}�<�/���һa�3�Y�qs4w����⇒4�>���n�i�	A���zv����ծf�?����Y���W�x�6ɢbs��&7�B�V��A�oĀ�������Ɵ�Q��u����$ã��;�Uh�%��T�!
is(,@|��M'���ß�酐��"�D��� �7�y�\�3���J!�&w����Qu��í���Wy�v��'�!�y%����#�̴�X��c����>��p�����^}Y#D)�]����	?eR^&^ff���N�����6G��'�Oo��î9$�Y���ݹ��8��;\-���[%��ݳ6H}���a��Z\�18�^.��D3�lDP���Cr���ZkiE�sm�n������+}�䉹��1�~��0�����92������ <˾�&������ -D�7k%Z��L�#�E�����w�Xo��0�Ω�
=k�q��_1j8���D��+f�v{5��5ٯ�{\( �4��7�/\9����8�l������_����(�"#ü��EH�ϸ�<�V=<%PB)}D��,�$q��x�[Tm�)�%�mb��%S�Grm�%w}"W�v��ҙ*a��惘DB4w�CN�|����bSf�Q��b|�1�:m�X�|��n���יU��A*�w�*ujT�<S���ZZ#���=tu��*e�7C��hR0�Nx�4��&��e]y�x�.�f�Xӌ�<V~2f����3�O�Z,��-ֶ���L�6r�~1�m�m�}��s�暓0�w��M���ɾ��,�@*��b�2c�@[l�>Y�`��g�'B��rX�Ȣ���)�����/��3����c����/�kY�m�5�{"�-��>�Rf&�U	��GA���2�^��c��E.dw2uqL�B���T�E��hN�_3��V�k����[�e��ڣ;��Н��&�ٝ8���Z��l�ަj��JqFxt_~�ְ �����#o��&�c���v[f����s���1J�+�X��Œ>�SGrrl�~G�u;�Ʃ���D0����cE*���B=ټ�����!�C�X,g#�pawC���fs�v�/�m˄��0�� !ם֩V����\�;�a;��67�§�;һ�^G���'�a�,����t��n(�}��ճfN��#�,\��Er�VT
Yf���d)��O2�d�VM,c@��;T�Qe�f)ə8�2@�IJ����۔�*�N��8�;6�ؽ�'e���.	}�Tx#'��?�b�c�mx�|Al�����,�	}��"Zى�x\`���O�9���`C����������F�=��5��� )
������:����N��4��fcw�>�;6��39��Xw�J�����2�yy��H>�
�v�?�f0�W���������g���]�����f��3_P�1t�+ d���	�dk0ʁlf����"�V�L��~5�{�Q�ߘ�̼c��.�
#�D�_ˉ@j~��^l��j�����'�儢�5��^��$��-uc\�g�r�]����Y����M������P�u.��Z�����{���-�4n�֝e�ٙWtN��\��杢�9*�]�ӣЧ���ۮ�ƹׂ�w{,8{5�"efHh؇Ң2��0ـS��ݹ$�n�^��Z�N�H��
_j��l�XTk9��[{qKA��R�&OfN�[<WL�޲���r�+�O�1j�j��S���9l���S�m�����D��:�ݿSu��`~�&'��=ͅ,m�l�DC��FqOn%YS7�[V��p��x]��1���>�;�jԗ�;����Ѥ6�1��kUz1���qqCJNH%ǚ��\GK�	�������\�A��^�ugM 	M�����e9�˖�=XPM-�x���2��n>�������:b�H��5���2��՘��Y(�xԟ��:T 9D�*z�mt��+i�X��\uI�� z��ǵ8S�L@�'�btfek}"���ev>���XQ��ؙ�'�.$vDe����d��%��GJ
<%�A{Ĉ�I=��s�c��Ow�A�9��U&/0��CL>�,Y/$,�\���<3ݮ.�u�����?� [ u�&]װ;g��;�-��*�-sQ^�$���W�oHƬ�3�q�A��.�y�_�cD��S̘�U� �Ͳ�"LT��26���j`����\��TT�n�}���W��g��F3�d�W���pT��l{����I�OOhwM@D=K/0'���)�0J�4P�S�W!}�K�)Q!f��NBvO��<M�u|;�z|�nb�B��v��ޠ�m��{�D���y���߿��h,��?��Ν\�սy��Rh�t|������,U�������S08~�[�1�ԯ͐���?�e�x��.�̼_�'B��H���j�話��wm��4�WoG�v~"<�Wt�r4j�e��wU�Wq���ew�֗��-t� ���	��Ӂx��o�'L�j����<�J���yIN���{^��n�h���qK�"E#�I#n�(��N�Yq��ZGE���¢W_��n�y6��&QXO�q ���O�����*#uZ3�^T���wG����b趖ჱҐ�%��/#.Z����{x#��pb����kƧ����ݼ&f웋�Ђ��ϖE��|������3!��'����_Ϳ��L�;C�Ԍ�1�=z��t��>��Q�eN��͢����g�*Zգ��1L�ϸ:'\o��/,��ll��b��DN\i�0Ox8��	�H�[[�3!=% ��#ѫ��^�-(�Fߜ�Cki�B�o��I�E����u��x�E62VN��%r��Au���u�;����L���2�3L�����r��TV$!�Ϻc����0O������{رp��v�ʭ/��M\�
���;�V��O$�Tm$��Y8af��t��h�'<"(�M B�M43u��d�`�Ma��R��j��w�<�u��G�=(I��셵?K_n@�v�;ʉ�W�D�j�|b�ݖ���.
j�:�A�S{�����N�o��q�q��*`��h����RJJ.A�u]�hB����z�f.d�s��ctl����z�3l��a����Փ���eO�'��d�@�Z��3
PT*A����f���e��:\z�$�DEAQ��WM�>�O<��Cfm�wU
Z����5��Jm~<3O�bt���$�N�o��6n��6��0��k'V⶯H�*��9XW�2��g�y��+&@�F�%�0�i�e-��R�]o�?��&вB�e`(M�m[*�w�p�涎=Nlfp���dt�.ݶ*��p���ԉ�ӆ�@:����4$��tL��R��!�q�,x���d��ڌ|�d:��`�5y29����5qq�5��!�Yd�7{�v	b+�K�|�v�c����FTZ�m�#a�4�/_�e� �/#�v����a�P�ѕ&t��l���J�K��!j���~���k�������5w����<�8��`��� �	!vyA��,�d�.�N�~=J~NS������dr��H̺b㥟��p�?��Z�|��{Qݕp�bRmbo�+����~��+�B�����M=��Q�.w��8�T�y��_b=�ۋTer;� yC��h!(V��f��qW�'��[K(R�"Y/g�8o!s�'5��Ѵ�(9<D�1ƞ�%��,g�Ɛ�F��~ff�K�z5�����S+��>�~J~��x�3���T���R<�Ee��G
5�n}
bo�.���nFq3
��[����<�c���&���a<(ry7Ztx��y���u�nl��-ѷͿ��
[���ʟ����-��4���̱%�T�*��%�f�y�(�$�/�a�u�]������Pza�#���~m���{�}vV�#��\�_x�:f)��f�L=�0e��nKD����|0�js:ٌ4p6C��ֆ�R-��^��Z�fyGQ���J���jf�F�kQxC�Aʓ�/�8F9Ue{l?��N�����`��_���;WM4D?+ׅ	d�,��2�=[�fr���� �U���~;ZE��%���)4?��V9��)��.1+w��8B�WHk���=��T��Ly
>Ez�N�r�F5�W�������H̥8�"L+�Y:z�Cjnxv��ȷ��1En̒K��r�+����2Y���ȫ��ayM��a�mwXޚM{�-�`b�`�c���2Эz?� �"���I/j�_�L+�u��f\�^�T�Y��������0�|W1$B�=�HA��6��TB��J"�١Ö@KI��	x�L���Ή������"��A��'t�W��2*v���IS�����K�߁A�]�b	\F���Q1��q���e{��8���:�'���c�x�g�� OZK�$�Pc�r3��2j�M�%Q�Nt�Ԑ���VO�^�j�Y!Vr�(@�7�5�����[f*���
�����������m��#�u)�̷-*��R\,� �-/a��h!6�jR.%�9��q�³gVC�b��[�za�]^=V��|��a���D7�~#)�v�>g.W��cl.��x�lCﲣ��k�<�1�J����i�G����/�{8�E�>�S�l\G�y�p�G�6�S��?:�����O��C?49��}��1�~�f$�AZ�c�{3U�r�iu|k��qc�(%=�5����v���S@�l�'��PK-Zk�#˳��fc�n��+�)�FN�I��:��3W�n�z����E��_�'Z�z	e���i^﫡L�N?��M��P3H�VRUM�؍�%Ǳe�r��+H�k�N��˰��#FO1���-�?���jo���}��:_�S�^���:xC�_Oج:�]�ٓ��g��r��,�N��^\ꞥDН��a����>�D�N�/Y��mG(�t���nnf_̧���堈6�娲�����F�U�ҞODVI	"=����W��NO7�t���;M&����l� �󁠤w���C*E�{8n�]��Gd��ΡWA]�zT���a����+6MCm5�8k.�W�?��_�~+���*���ǆw��J�������\'?�":�fz՚�pv�*5���#�FZ	�.a��4	��gR��v3	+���t�}\�st$U0�>nWC��NR��ݶ��(��Y`3H��&�Q~��P�q��C�]+<6� j���3�#�Ez�'����#����~>�=ȃ]�ż]lB΃@f���<0��ք����K�C�W�<+�_v�b�ؠ(e� �Vt�0�_"]"�߅}-�[�[l��zڱR��IG�m���H�Mqï���Ս�I=���K�W�1�fF2R���-E�p�g�Q���xP�ɘ����Vɇ1���3�on�s�������g{�p:������pe�`#]�p�������DT]��)2���L��WQnE���w�Hc.
֕� J
�ftn�º+|6���� e^��qX�9lq6����F.�Ojh>�I�KU[��u�h���ӭ��ۄ�g��q�Q����Λ-= m@�eη�\j��w#�C��nTx��>��T!��Pԛ�Y6��_RD����^�bH�p_�7�1�O���(��q������_�H������\Ō�Fz`~+z�Y�֔�ȣ���-@���*��]q~���<����߭4j�m�w�Q���V��pr�S���߃�� ��<�i�Y3k�='L�X$d�{o�Dy�݈5���cI dmȷq�2J��"_&�P��@1.T���[f�ܵ�������a�G/�M�BZ�C�q/�r��,��[�qyǂf�*77;��{�`�tH.��`ڧŃϓ���_�8�P�zY�B'�6J��5��M�J�A�^Oʋ������(�G���J�Nt����k��U��V�����(w6�Պ�z�w5SQ��h�I�hV��1�p�d~7;�<�_�du7�+ �,������uI�?�z����������Yt�c"l"'WS�ϝ8H5늘�	���HN6x���dV������-�{� {�pv6%����8kt�p7� e5�W��?��z�
�������v�������P��2�2[�TA92��r!�p8ć
G>���#=��_������OZ��}��~)l?;��|y����a���u����(�q��K�ȵ/��,A� ߙve�'@E�{dۿ��4��&4��SSM���ZZ^�w!%WL�;������؝" u�$�H9����햘;�
�!4�eȚ�3S!?�<t�ti8IF����`]:�>	�3��ǖ7l�f�t\��4��~��N����w�r��c����_�x#u�_����ɳZ��I��b��ꄖ���vba%�Xk�����tu�J	�-�h�٬ow�7j���o�qCah����)�H�<�]�Ш~oCU�z�9�o�$TQ���C�;�\�(L��%�ǖ񏤽�i7� _~�_��y�R�cW(�b4�x�;<��� �:�����=��Tk�>� ��/�F�wh��[��6�81��+�5X�H�h�u�I�Ѻ�So����Yg����V��!VkK��)��~��� ?�ƣ~�� :���%��>%-�+�P�-a���0��	��G���J��_�SG��l����'0~�R]�(u@m��9{��EN<���������؝���ME������Y�Cm�_HB���"V�I)����_,����<�lR`c�P�~KW���H�*$*�f��_� �+�{NqWJb���xf*�����y6~�)��i��`AЅ���\y�"zQ�# \#�,I��Wچ�Ӯ�����&�Rq�˼K�oU��Z����:oFZ��\�@�|-�k�b�`��MtFE��Y�K���Oriƿ�o;�G	NN5�y|*Y��/�p���7EF�	�Ǟ�=�$~�lYBm�_�\G2
�p�<�mnϮ,����St|6�s*@k�����{�Wbw��[F�Z7\�L�*�^PNg��.���F�� �E�:�e��A���2z�D�di� ��a���rlde�:�J#��h���"Zcy���P*�4Bi@f�����J?���Ķ�bBCw4�G��/���f�6ڧ���$/�N�J���Y$K�Ѥ1�_��O�U��;ן�k�e�����iD�|E��J�BJ���*�����[�T����>u�ii�0xmR��A=܁��<����s?4�TA��D����c�X�Q[xr�VUl�h��"��]?k�kM�aC
�}(�V�J=̚(^]�/$�R����C�6�Ԛ/Q��i��Y��{Є�!���ΊC1:9H�>�����!l���n����Q�<\:���)����*�U�+�����������6&ix��9(����qC+L�΍�Uc@8s%�T2v0�7�A˩���̹����`��*V��Л+��VT����^���0��.٘��,0�P�4F��q�ИF���O��S\�/ږ��L8�V�Q�9�/� .���rnqo��
T��e1	"��Y��_<�n#�[k]�>.��>vV�'���O� ��&���-j�|�Ρ��5� �@�Re!�z��+`�*[7� (�ӄ�Uۏ����JrۆL�@�oR�}��P���#�_��Qб|�X @�>�;$uW�¶\�&uw�0�q��9��\]N�K�⎸�A����87����� �X� ����z�t��zS�D�k�F��_�PNe
i�g�e^{]�Aʽ��0,:�|�ʌ���3�h_v��]�ê���6Sd�)�̵.�P�y���sIy�\�1�x����A`�a���!���>'��4r
bЖ��>S-�}��H#��ز�z^�?^\���q����C����o�}m��ʃ�џ�.��W�[[��,Z ����V�p�+������Қϗ�Z]W�=�,��_��:>�v��0c��q�SL,��G�q��5�YdE�O�����|F�D7n~�P�5�W5R���=�9 ��G��+Ud�LT�? �{xp�q����HQ�m���{-�`���s/���SJ�}E����g����>���,�7Ԥץr��#4�-�����|�j���sL���GO��f����󸨭f��f����ك��ґ�JM���vs���ʜ4�Cf5��Kп�"�)���@��i�*��(;"[�(�S*��L7�ۋ��.����e���@��e�y�� �^��hU`"�1�����	&�&ڣ����/�Fq��M�)�׺��ҥ�ʉ�;����om}ǆ�e̓���j�ϴ�G�����2���x��k��L�-���T6� �����<O-�|lYr�+�'��9�]�R� `���Bf�*��!ߣ?��
�wy��{&&d���\���o�Yp���bFֵ4�)����zs9�a��Ȋ {�c@�{m�~4�,�{!�ρ�g��x��A�8���ep����'swyr�&E����-�@�[J��B�^�V5p����5	���UB��G�!7\�]��5ֳ�|�@�GY�J9�y@�K�1^<I~�y��36qSS���%Wb3� �� "�1Dn�����ח��J��D�w���^'�N!ڢg�K�k�&7e��o�풫��9���)�R! ���{�E�yQ���Si�='6��i[tͼ��H��K@��K�m?rEma��}'��,/G@�࿖�p��N{�<���i�SX+({I]��3�s�H��e��G�/f�W���H���xN��y�G�^D��Pv�z��$}#������h"����j���c �8:����k���Z��|�]@=��K����%�����`��N�/~(O�Qt�3�R�Yo[\ʲ�![�B��:��d�83�Y�4��T���LZ�et���@����� 2��kw�oq�0,J���g	�0��u0�0���^�i�˂�*,����+���H��4	��ACz�v��X�ir�?�?��ȓ�F`|H�g��?�{q�{��G�b��;E7�^m���:����G�
�4�/(ؑwN�f�^�f�w��cU����y�ds��G7���ݏtԞ�N���WSi�p�z�r'��J���t�+?7��M{�#��h�ս��s��`���=r���z-H+Q�2b�~p�*��{�����L�?w��.q��.g1�A
���p��*['�]ȓ>`}�.&��7
��@2��4���8����쯐���#����M��z{qhI��Q��lL��"B3����t��:�ʝ�G�
Ƈ�-���LF��kDq���lD`SiA��f���~��������;��}�лY��zj���^�%:��F����z6fBV�ٜ��t%�W�[����	� ������J�!b�/���������6m!���N�=� �� �{^&�v��� d��QP���%�	Ɠ��%o�ςS
��؝�����������JK�edyY�GZ�j�XiS'v�̣p<��=����>�tA�'��a��E@�~ځy��4���>a)���b��+vB���p��3�T�W��E��Wm��:6p�n�+�t1'Ux����"�����&#��9���v�ٕ?3���N<)� 6j�)��?�-�o�
��|��N[�G�����!��4�D'OS�"�t1�{�D�S��Ʃ�B](�xf�г�X����H�q���\/��m��D|#╉ޖ����N6��`�!�.>�/c�S4+D���RXA���;ςYd�7��X�a��_;�=�h�3�[)a���_%F;k�fL5���j���;�~i1_������<�=��#����gv����/$�@q���κN��@f�63_g��L�@��|����C�.��IX�n7��蔢��j�t�h��`<�!����������՜�;�.��x�2
�0��\h�c*�zw�h���p��\b)�~q��4�z����VW�^���ȅ��'m�MF�{�hi^��b?J��ڝ�u@�w��3�}}0��	3�T�m�g�ڨ�֞8�p�3z;�����xS8Y��2�w��0�a�oN����p�Ei�����Y����ɨ�1�e`��m�>"ec���}52��_�\�z�Pu(/�Uک=Q�o��]$H�Gw�s}�x9��<�I�j�w6��犢�Gp�3T����.��㹘���EZ4]gY�� :d2�{��j�n�~������޵v�;��@����.�ğ�S8d+/I"�Q	R�C�!��w���H���CX���f�^��ۏ��+�vI�3�ND+��t�kj�N\3Y�K�����v��0�/i�4����AK���8H-�d��@���Y�e�g�]m�m9��б��D�?S�M�<�
u�~�a��H���<�R
5׾��i�C�褵R�*��F�n��3e������r��Dۗ�R�ʐY�*�}>�)}jL��S��Y���Ԡ�@w���u��'�-OR͛2�H��@n����(f�d�L fƫ�5C,qN��5�ng<�W�*1 ��L٬�'/��-�ႇ6`���j���������Z�&�!~�~H�C/��x���w˞e͈{����/%�>͠�OzY!���R#CЎ.2�{�5b���J�9�X�ny�b��.�eu1��M��~-e4<j7W	e�i�[oK"T���P@��ý�X�r!��nM�h9�����KY��?��L�f�CKߛ�z;��������[ߦ�J���Fr���.�z�	����m=�#��v���Ȍ�m����k���y1����9u��V ���zr�-�G�tג�X�Vʍ�0�A����]��^�
)�?�蕧[�_hVwH/���
..4,��ڳ�A��{iz!۩�Gz�![Ť��c����{k�`a�M�hZy�t�<nu(d�UC�����p}�g�ُݵ�'�ζ���z���9v́w_��R3�]�$�Pj��3�������пR��{@Rz0��E�����xb�ӎ��y:S��j��% -[_Թ�ޗ�UBu1�y�t$�ݷ���� ��z<<5v(ǛN�f�ڔ����O���z�Z���P��uO��M˃�L��ol\	S��z��f�����[N2ʫ�����J�R�U��y������- <S��/�a�153qH=��v{�ͶBݦ��j-��	 ��b�&#EX�R���T����'�O�*�y
�W��g�	�y�\X[�|�(ң~FIUYF�9"M%s6%���KT��W�*�
`��-
�%��lci�X�܌���:��C1]|z�����J�$`��W�]8S�vkx��Z�s���u��$Y�(`+I�!�����T��1C��f�"Q�Fu^�6�Y.��y3�1� ����Ol����HZA֫(�D	�d�L�%��p�f���$�\�]��[V�W ��+6�&&4��+@1~�Z��z-O{>@p�s��VK�v����y@�_��zַ���6B&��TV��焔��Ho{�G��%JU`Uٰ� �̙^n�(�-�s��/]�J)����=�Oq}��A��7�<3�8��rO�HaPް��&�H #zM�Ғ�%1����c�e�=ڋr���x �^�a�w�ә��j�`3�N��PK����0�{K�E����"�(�F|��t	��λ������,�H����"�&KeI�%��`�Ab'�xdL=Su�V�G	4B����:i����GIU0��-�W'Ҵ�SQ&��
hֽNhF�J�@�;��ktR��k$�����Z�0~n���36����sB���Һ&Cz��t�i_U�h�\Ph���A�C`�<�V�Ԇ��{�l�qM21�~n�Dn"h 7���6x�i�NШ����a�$3?����H\�	Q���$=Q Y�A'%��h��u�h���{7K�8Ԓ� ��T\��S3���r����� �gÊ ���U:�����}�i�$�Bl��{���ֽ2z�
vA(�6��/w����E5v#�չ#E�����Hu�K�H�"_ix���[_6�nN1���6PU;e$1�z0!��x�9��$��b��}�/�m�n��/�M�<
��Q���B��ϝ�}X���i�\r�^���V?�7pJ��5x&���F?��ʘk����W�j�/��߉lH�a_L 2a����>m��*1�jN�m~��z5���;��0o����ԍ�o
[��;�*��#�Y��a�o�"/�����oQ_�i"�x:GRGf��V�����4���ɒh��zc�A㺎�����ڣ��f�ߎv�y���~Ot��]�:(YE�D�9�AZ����ᾡ�?������q+01SRd�L���}�N j��ro2��^�G�qX����]�z�1czŻ�Ti��Zr��F���vF8~�/�5F�cJXF�E�1`��4F��<�{�06 �e��E�O�&��o�ɢ`��ř(|�GV=�@���+������P�)
ڹTtL�X��^+IU�裷�ĥ� -Q�m%^�����P3���~	QO0G�h��~��N��9u>9����e*sc��f�H��[\LZ1�$*Ze){k���&��W��8㤚"y� �0��h�)�H:�cV�DP���4�.���w��x;�=��]����=x;��RA�?�i���;8�!fp�������'M
4F�/.�i{�+�����T/�I�� ���7��Ց]���kc�w�;���?i�\M�5�W՞������q�����f�=�X��nV+j�1�F+�d�B��Jco����9�����v�vx���2��� Q�`��=V���ܻ�5�G[9���b�ƀ����p��9��a@ּ( =���v�e/��l��6rZ��4%��J�3JK��V�A�Am�RV��S�ɇ�˜���a��g[���_]�6�f^��|�b�a:���v/�`=�c&J.��9SC}����(q/�6�ꠜ�R����a.D]C܄d���c��I�8R9�P���Pl/������C���@��.��[���H6�$ݲ2������%H_0,�Ŏ��GɉxY"�w
��9�@�s�j�k�C����̘����>z*ūξ,��y��j�G�ι1���]}[ߺp����s3�v��t���^���������w�ؖ���NN��'(|^��<p˃�f��F)�т�+l���)r�
c�����6���Ț���[+�y�J�m�\i�����]Wf�M�ׂ��vJ�(%V��{�Vrs�M� ��v��dm�m�0*+w¨���ˤ�����8H�����Ҟ~f��7Y�Ǐk�����^��-Rފ��%�VhJ�v�{�{\N+K��1��_Jv����p� ���Q�c[�toA#z�b{d$�wi�>�Y����z�.�G�3:zil���O��X+�&�Rtu����Py5��E��F���4���ww��}��K�X�z�щ��O~��d�R�rY5)�>�A_W�����R�Y��<�a�E��:Y��zsuh�şl,q�`I����T���b�7�ʖ�=���A��n+� �h{����>B�푄�y����*r�_�
��Es�F���^����y��ɺ7-��>[�Q���Յ�]&�f����6�ѽ��̄�Pf¨������S��d.���,i�j����f$��A�<�6'v�*�㇢v��D�F���)aV$C��&���QqV+���_R�:j.hyN)h9C�=��W|�����Q�U�	���W@�璞ROe�J���X�����+{���ґ��_p���\�1�̝�W9�
+Ujp�.�����9�1��;ڵ�ԁKu���y�o93�Y7��:ܘ�<W}�Ē(+��n�Å�wIl���OE�Vi�^�b|������ܜ�Įy��΍N���A�_Tk�*����bV�R��Ƒ&H�bɗ1屒�1ԉ�#��d�i�W����xmף�(��I�]ܖ6t�s%���T[�h�U�����[|�����ֶ���c����ɛ��~A��hVt�\�er3hl%�LK@��e'��;�P%���C5�@��p�x��'��;�]7*����X�$u�����/3��˦��~�t���y�m(��l��d�H%�M1�k"#�+�o��f1c�Ƒ\�1L�|.��Ws��]j'�K��"�u��{<30�8_���;��z�ݮ����q�"8���QT�K�>�)S�a랆�̾�~ZM�0lTi�AC3�$���\�Q�seWK�L+���ԙ�e�Ɏ��96}�!�ڐ?�F��{$���~��@�(Q{��z>�ꮊ��f���?d���x(�\����F��fdg�)��9�RF�z�mv��5�d��c+��1%x	�}����2������^�S<��?=/-��K_Mk����Ύ���M�z���V`|zBZbxse��ٗW��^ҷ&T���HĉW
[��[,xTG��0�:��!_]�Ç��WDU�UN��@Ȋ�P��>���z!��z�b[�l��� "����v~^��z���0	�ʤ���ƺ�ݻܺ��Uߡ`cc�\n���/�Nr�z�o%Œp�h�Ou<��w��w�>씽R�͗�r�lw�D~�HT�
�!F=>q������N/5&����+��`1�Ȋ���V�Ni9(է���2L�v�f{���;�����q���
RGP�bA�"(]Z("�CB�0"HS� �I�t��PBI��@����n��������keɊ����g�}�{��t��d�j枣�i�V����&��O�\���+��+D�C��,��^ee/�Ra ��>D�I)ڌ����D��/R�lqr6�\����[����&ꚶ�Z�a��V�� ��و{%=�b��Z�'Gz#ON\�s+c���UyC��w7#e����baE����P�N��_�ߡ|3l��E��:NBmH�7���:���/�?z�{<J��k=�yw]܍9y�P�,J�5���?P�'��3 �i^��{��Si���9{X�@S+�4k��t�Fڑ�/������lEQ��������cIeQZ���*�\��Q�v\�x��
q�^!���;j�yz<8o�"��N>S(��r�|E�m�C�����J�X1�����e� �ܥ�4G_�w7s۩kG�F%H)pW�j�ޮ����&��>�x��J(�li�?��?Í�)����!��L[o.r�yG�����.�&������I������5���K��y�|��?a�.����몘q1J`��M�J�n>Ӳ�Q��B�Qm���G���d/�Q�(�!1i�O�X⢒/�s��VQ��E��K�(����/��X$��g���]}x��V�og�kF/���]>�P��u]n��W��P�� ��f���qn?u�>�.j�ʹ��(3�8)I����'��� @���XD/5[f�e���W+Jt�cJL.��W������䣸��O�xY��ᦥ��a.�y��P��Z���\k��J�>[���!{y�r��EU���s�u�~���u?[T��,
�Q�*��ل��h�����9�nϚJqf`��P0��>�!��@���9C�>H9�`V����)��4V4猤w�uF�Ĭ��<X��D]�U��vs<���7�GA��*�}r�C'�����c�%�4��C5��ӱ�=�se��.j�I�e�PS��!z�RF�t���,Hg�i96�W������i�$�Ѷ���:^����XdGh��=v��"���w��t�K�ш2��T�)1
Y��F���{�ܼ��H��3��
�Q�1��}���`�k�u�|��4B���"�K����L�N���<�ȁZn��f�pD�;U��õ�-�!:��Vݗh��?pr�ߟ�Y\�$*���w>P*���NQ�1�_��1�q촁�)DD�p�6��<=^o�`�:���@���ݿ-����`|Z�fG���s:�4��� �i+q�,��S��V�!}Z�����}h�i4�x�&�l��K`�^�5.tH��ѡ��}���k_tb^���;�y��ie��8NL:�wL6(��֍��ҀTs��R<F��.#iN����X���q8+���������w��i��?��*�[�}PR��q��g�������
���̃zs�'��Z4�z�w�_�@H!je���A	e�J�탇��ɻ��G�L����S�1��Z���$'3f���L	-��9��c#�����n��.z4f�q�G��6�����"c?5đ7�5��Ke�;ṉ����u��U�Z5�H��27�9���,�����J��@������J����×y�xL�����]���vr,�.{cR��渂��ī �^�tP6�	��KY��὇�	`f�h�(�f�[s��M]�yFy�f�V��"z�$ZS�^e2Ҏ�����2>y�0�Z�ir�x�n|�]�}��#���sg3��둲�Ϊ�!K�����MZ�)�1f�[R{is�IPCPw6���J����f���!���<I�ؙ��GƇg�? p�q>��_kt�\<��]L��q�~s}B��KİF�ȱ��������F=���K)�ŏ�l����p����u��vW����R�?���3fGn�i��S��G���ڵ����|� S�*�P��A��U�~��D�l-"�d��� 
S�X��~�_���pN�������2J_��;Q4H�u�W�/��}�<�kP��N���kd�Ol�Q�m�\X�.�b�x�����͵7Fܗ��)����,dʹ����X9�%ݗ$�c���v����Y�����`�wJDw��;*���S��3'��
���d��Eg����߄g�|�b6侣�!���'W���8��A&]���##�4k��ٟ��6.Au��H����l[���+�<�@�Q����^��F(Ezb��^��d3�X
D��7i�!�7�+M��'��/y��B)>�z�<1j,��p�A5�p�I)���勿�����[u�u��BϏ׸�\� �Zף�����8ZWv&�'�g_w=3�?�����B�tu+@ �����2��U�ox3S=���d �4��0��=�2m͐Z�V���嵲)�1��t��.>����ס�Q�܍��������N�,�⏦n�S%��(Z�����Vv/za3�����q~2�I��J{�9"8�`I�0z�[r�}e*��R�f��'�'/a�o~�i��z\�\��tM꽪�\s�x�h�� ����2Pk�K+�K1�ܞЬ)�Va�Prk�k�]#��	��Y�)i�$�jJ������`�i��J�c�^"�8����זi]��I�la�T~w���н/`�W�f����U�^��� �7�׽/� &7��I���i�^V���k�U��m�j��!6i����71�?�5�Ѿ�W,��i��8��Nm�ں�w9;ưA����������[ d>{�c�5��8�m0�A��Kz�'�����tլ/sqG�J}�n���@��m�ɣ�C��ۇ��؛�_u�Wd|.]z��=$Ӕ-��q�r�%Π� �z�8ݒF�[��I��uh���V��	�q(+��;e�hȈ�:d�:��wI3��g	ʷ_u�[)C��a�"�v�s,G? !_���z���9�^�zUL���.����O^�0`�l��ܞ� \�BX:��̬�ѠO�h�ͲI��eR��p�5R�DU�	�d���:��#SNC�����,q�*?f:\c���n��w����_<�Zd���] �Ru�@�ߺ�ӵ�������r�>13��Ǯ@����p���њ���N�'��b����z���'�����i�JP.��̨����5;��H�I}P�����{�Jځ���t-�ı��3tM���]�;���F
r��ݍ �.ǘ�uՉ�D�"��s�c^3kO��6���a:�n�>(�9�JR�t���N�Q%U��Co�h*����n�Lrܨ���@�K��3�X����ҫ��<�;���}�%�S�$�������]!�/���}D�b�j�e�+�Q]Om4ǟl�O��0�?b�����س�49�\�l�ޒ�?\]���:��������ջ��^oVn4+`�B����ȷ��z�Xc��_�K
�K��^����f�j�X,ME`��%��	�:�)q����4mᵧ��G�����W~�՛���"\jZ�����o,9��*��`S߆
�Mf"F��O�b������zL��ͨ�*���/��]���Wb��}�W%V���, �ߕX9�) ���A9�K�N5�ĵ�O�a�ٌC�51,�Z���1%JZb;F-��S��	�˼�� GF�\��g9�|����ËΜY:�y=L/�6�{?�\��=~�������<ﭜvñ���
ïUU��~u��*�NT���ri;������/b������P���ZV� � �[�O��>jN;�P�Ȕ2�����(#/�o�$q`{3|o�#26 >��ma�	N%���Y�(䫋�ah@�c�+V�\�gb�����o�_��j��?~T��	����?�/�6�6�]�o���9���@yo�oh��CQ�G�@lt8��ȑ���A���ʹ�Ъ��X�`:��9�}W(+�Q��$�>������ͱ!�:�6`<���e���_i��s�?ڀ}�@�|�$�?jF��V䮑����,����S)���r�?��Jw'��U�U����Q���8W�N��&�X�G�ư��m��C}*#�K8�ssV����jUf���fc�a�-!�Ce�;DGJ"Y'vW���.�rhX�������^���?��A	�{A�厾T�
�O�����u��όK.%��<)!��yZG,b�h��у�����f!\hZҖ+ХV��(�h�w�"c�M_�aw}�CUT	�2���F_Z�.��ӌƽ�yČCE��R�w�"�_vm��'��g>��E�/�}�o<��Y�A�!����Z�/?��hf�`�:�<���| ���Ŕ<�iоC_S����OT0 9[�����Ip�\��*˹a@��� \@k(�{|:�:	ޢ� ��۰��{�=��dasQO�~	����p��0+��P�22��5�7@��g���{������O� �^�Zyp��0��L���?�,#��*?� e�S�,sW"[�,9Rf{�=d]����u'��fݿQz��l������p){>e�X˥6o�E',i�6��(XL-�W#�x���zŔ�P}�]�6(�޳}�n���W4o2��\��ֺH��WRc��m��$ ���Q
MK2�%|\8eտQ�}�)Q1���zԵ�2�>�8��j��z��^1}�����2�eʹ�7�.�qڟ��M���dյm��� u�)�����a�M�������=����_7�b+JWh�:���r�W�uP���7U�w����� CUV�� WTu�愈w����	���ܟ�N^t��c����s_�P{1I��~�_���<)i��6�7ȧ�{��h)�x�U/5���?�������1w�����n�߭������������֓l�O�C�K�Y�:�!
ލ3�zqzEg1^	�������x/ �v���x��g��f���N�{+3M��vj��d��o3ٲ1�W8��ǆ�$+[O\�/G���2NW��\UK>ET��C7���?2?��0,l���Ľ�8�w�(*Ų��vW��5�W��M�/�¢~�ňdۧ��D�o��$�G[&=̔��h!�-1o;ۗ����aˮ��&�k��Qs{�V�`�O��p��Ɵ������;��#�9����t�����W@�/��owH~�p�x��5��%v%�3zg���A�6Q�SZ&t�����qWY�[9��W��Ų���B.ގ==n�������)L:&��Q�����h�z»�h;Qּ�����;W�a��m�QD�T������S,֦f�����%(ne�*?��a��D�\�my@2Y��\#�,�lu�������jWŐM��#����H�����D~wy�A�$���FW�_�(j�`ߝ���@ݐez���Z�kx�\ڌ�8�Q��h�\��E���7���92�6:��)����������9E���P���Ĥ��\�geAtX����i�������ZnƠr���`���g_KI�3�t�3�ҁ��]dr��ޠ���y��]��H,9oL|Y���|��|�e9��"'1Dw;�;�8��G(%W���=��v��i�*c;P�h�I�\`y�ܬ��s�gl۞"���ִ��HO��~��ޜ���YU����Z1c�g�瘲�����D$��]�Z�b
�b�~��t�Q�d�B���f(��HC��xGQ���	���F���\�@?76_^��?��>N�q�Kg��m,Ҷ� �<"�R}������o����gP��F�R�ҡ�����꣭m���R�Wá���\���0ky�H��V��e Lw�ri9�)��c�3 �-�����)��W&.J/�s�g<�����Ыls��<�1\j2U�� ��ņ�7�����N�N����QwHoC?��zC4o]�:�zk�=�<zGٙ�q�zo�}��Ϸ*^~������KtGb�&����v�Edh�%N^5��U�k4��M�Z����������f���)Bm�	��O֙"}U%�b�2��k�ş���Q��h��lu�+=5�c*��@�T�'�2C}��J���B���9F�AHZ��̈́�_�=��{�P���m-g������EHL/����5�Ǻv b3 ��Ss�vg��|� ��k|ʛ��N��W��a>�J���c����p҅��VS,ϵtEx鞻2��V�_M�{����}���9h:��ל��m�%{�WЇ�
$��:��K��8�@�#>6Zn�w���z2��'�܍�5��3ф�EE�[�nI��6{J�7�_o�<��-����T��j�����jr~uy�;�૒*�$I:�O���E��}�TI`�_/{HS��p���2�������K?����I�����a�?N���;	�7�����������@G-b z%��D��G�p�Kwg��$D&��_ ���7s �@	.�C7��[w�/wQT���w �FA�Yo^WۏY�r�d�C���U���S}o<A�uD��ZB���g����!T9`I�IR Dz�|>�����[�h�*2[���ϙ���*�o��e34�YQ�)�.", �Xx6�*8���쪚"��K7= �<M�����%6�E��y(x���rկ��Ϩ��J*ו��t	|kJ�P��2��֒ɪ�QTdÜ_�ͪ�X��=�1j�2cC���QXS�����?@X�qEOI��j0�|Y�W��Ԍ�q�Q�S���:f.���Η�'v�[늬4��Us9(Hp���%uЯ�-�\��s	�S8e#>�	t�_}Gn-�gQ����M�b�|Pw��b�@�����n���T���#��d��J9PG4����e����0�G?P��j�X�'�Ĉ��x�i�}��(+{����3�xi�-g;�^�`<��q��P�?�F�V]�,�^&ל�œ����\
�FJ��MO�ߔ�u�u���z�?���ܷ?]�AYxv*��l�u�S�x���2W��E��r/[�d &������Uwj1k��@�:r��#��$�������¶䭭ETz���̓���k ���gi_��~�U1[�Y��J&$��Xi]U#6��
��͆xw2�Z�^��)r��"�N�=�Պl�����X����嬩�t�H���V2�,�޽��f38�Z�0�R{hX�7&?��;�����lFD�W��J :���b6m��4��R�a#��=ee����ѧ�.�h����I�C�} ]M&�p~���74�G\7��|5��n�� B\j�PSESp�>�A_�_� ��R���pֽ��ՐGa���W���$$��2"K��n��.�����K��'9���APa���9w�2&�d��-����Ɖ˧zoh�$R�����&V�pKbR�E��l~<F|�� ���N5���UHH{#��#`���q���XOm�:�V����Z��not�Q�Q�̀���!�ŲKq�����j�T�0�E���Wr��*!o�z��/;}� 1{���u��#:��s�L$tO�֨aN��?����=������Q	�[˛�&�����n��u�'�I�m=�)�Y�K���3#&F�댈X��Ӎ\�-��^��uC�̙�:iRz��8�%p��30��ev�~2��G�J{g���y��_�s\6I�t�s���_0?��ڤ�F!#��r��Q��Ɠ^��#��sk��(�����}u�� �-Ǡk�5�tE�pB��7Yf/'o6dvH2�����i�]M�uJ��P�)���`:-�nꭽZ��wT����URo���MT���g��f�=Z�.1�|~~���nq�b��Y��g��
���'2s�s�r�o���&��䜹�#@8h��ܺ�Y!��J���K���3���`*V7��}^�o;'�5�RY����N���Х�:o�Nѵ��e[�����R,R����w]?4k�q���O����_��\;��"q��5�߇�z�}qJ�Ѐm3��t	/c�Ύ��hG*e�g{�T��2A��7��')E�l����F��ҴkY��4����T?l
�q���^��#���6�t��Kw���s���ً)	\��J���ye������A����(H������d@벇㞿y���9|g�y�!V�z\;}s��"Z�'�_�|���_�d��S�,�	���&M����y�D]���W�/��M&N�#�fZZ���R��Ͻ����SJ0��m��}|�_���$�6�*�W��rC-�$v�r��A��Eq�>Cp�`�����K�T
Rn��~�a�3�=H7����O(Ÿ���rk�f2||<�T���� ��!z��a� �3�_�$8�s��$i�tӧ�D�hx� �u�A?�'���a�ㅃ��W����f�%ۋJӞB"��^�3��M��:��\|�U!�F	Y��)h?�l��3�3���%M.s�Ik	����0��8��U]�^`&aZ*�{�cqi&�A�n[�����qy�J-#n&܌�@e�v1�&���#�W���1����k�Яj�6��1��KS1��*`�=��gZ�B�H���ؙ@��f�;��2�e�U�y�߀#l��y|g�n//��\'IJ��v�?fu
���+�ҷ�Ƨ�wė8D�"������q��/v� �f@����� on�����A��R
�l�oR�o�0G�-�S���B��!����y�XIm|���<�i��͕4�R����U#m� ۥP��♚6o�R*���è�̆`�M���qބ�/.�����=��Y�x�\K
�>c��������E���p�n]����B�������u�ܗ�������O��Yc/�� H]��}(�F��o%cDW��珿\&-����6R��0�S�2^�鹙�f���&���E�-m t}��N��N�ė5M�؄�Q����_Wl�������N��2��T+}�ڡ.IH~�h�n�/'R�` ����oh�%��Q�L/�Vl�T�h��Q��x�ВG]�.���bLm�^��m�>Y77[�o�V��C¦�3�����'`����m�A B��՚5�(�]��'k'" �p��w��N@MY#�V��%�Ϡ�N��T N�
)�qX_АL��p�>;H�4q�+6���������4V����^3����o�2��4�&���EƸkU���)3$��ӋM�P�~�@���'����\h:lPR����t�]x=qn\!�( �+������@~w�{F��L����t=r��6TH�#D�Fٳjy��͍"L̥�����Ӱ����;n`� ���t�e�+Mޓ� �W3z����\�A~�5�mVW.�l����3w�03��O��������N�DYF��ƕ 5��'�����ڨWx�]�E�Si5��~f0�e�����&fN۸�n'Ћ�9���������z��i������`*�ST��S7厧�Ⱦ�U	t�i||���.*�\~U�65����i��DH�|Y�����׏S���,Ges�ёV΁�?#�H���Mwe]�&�r:�����A��4Q��,kܜF�#�'�y!^a�ѓ.A���l�u �qW1�JS�!��o�'q��ߚԯ�8����:��$���a�����u3c���4x�����M�_�6��Y�?�SY�x�Ϡ�����"��|��-�ʍ1?��k�{�2U�ݛ�ԉNNx����m��\�e��4���T�B��n�:H��W�6�x��W~q�
�Vn�LgF@�:�u)k9�jb�&?�����6N��yip��͙E�Y�J��bʊ¦�~��� ��/��1Z`X�"�F�6�d��,��
�|�fD��Ju��gԂY��UԿ��[4!�J�Y3J�����0⽚r�y��w=��H�quW�[�����~�П||�A�!��LYR�� �0S �D�*�4��+z5}{><kGU8ڗ���H��Qܬ�Ui&� aE[��0TG����J�MB3l�_�2��Z��(5��A� '|�*IP��YnH��h(���F�����,����u�+]3';i���BO��@=xh��>���	6�����1���g�Rt'�}t�S[��i���V0�zEF�ɟ���R,�k�r�%����dY�B��}3���."�;�4h&j./6����R����Ƕd����X���/�>�����$���',�|+�vu�U�gE,u�ƿ��?�����O�p�T�;�)������c�^��v������|68r^i����Gz�tT�l��	�'�7��>ր��D{�.�y��vhy��*����s,/i!��S�Ȓ~/P{ݝ�f��m/�Ww���6�B�z�u���g/ڡO��N�M��θji`�%���j�r� ��sv��k�)MwV��x�,��7�s�;@�5i�^�)�K�|C�# ���{O�r_K��?��0ܿ���^�¥��#��#3r|���EO�c/▹q%���p�1y3�!�_E
���������g�WvB���,�#l>1& �,�de� �Pm�"��h���+i l�3�,��B��3��&�vb��]o�=�'/�o�\4����*TX�y�K��B:ɏ��'ԯ���M&�5��(�U�{�Ŷ��G�rz�|� ���V���4^8:Q{����dչ��b!(�B~�r+������5^*O���~��ɤ�V8g	��n���	R����cy��nM��������^�ϥ/,N��6L/W��U+>�s��Uf�S��\Ƹϯ���ۚ`/?9o�<u�r�.�K��Rf%q�hm�$=��q^�L[=)%K�$���K�|?֟Zu�8�K��kL�C��[T�� H��kS��'Ҋ�K��?�0"�.�w�̾��+S��DN(}~�g���'�H�B����S5
�};�M�������/F$sҎdX�Ed�]F�iQ���sJ����,e��]U��9��;J����]��R�O�D9��{A{EU��y�p)�{��Z	
�(``�� ƽ��O���^�YX0�_N6�QC�LB:%k���\��T� #�%�G��u�4�&���i�VL'q���>2��Ksfkg��>{��[��@��f�������E�JbQ��W�>
��4H��3%���)$D��0�Tt�p�tN�o�%����%MD�a��C���=�A�(7Z�����u��:�"	R<H�Y|Ë�R!����'b4��U��̍ˏN�|�B�˖_��Mp�.C����H8%��&GG��{�3��V��EI��5�q�OV>-[�-)J�d>V��XE�F�V*n��6��+}9��,EL�Tfi�g�3�������y%��y�������0�*�pR�^��<~���ک��9�/B&u�{0mo���K[~�����Z�%�2�C���)��ű�Y��Z�˪�
).���A�F��^��;_ά���:�$L�����E��둯/��{5�E��`X�z�R�@<6��0H��z�k��]q�V�b�J'���n��nU�\��0g,�i�&����Wd�l�V�F-��(�|�뮲���l���	���ݼ;����&1�ġ���n����9�����r�X����#ې%���@�=}���n�:�vD����?H'�/�6G,����p�F�n�F�����N6 �@���_���Z/%\�D��q�y��� �÷���y��5	���F��p�=�Ҷ����U��ϯ8k B�M��G"��H�Ź���3�\;Lw{��6��VW�DR1]u!�*K�;>�[������i���gF�^��LϺ*l�y��B��:����������
J� ��=��H:��'9�Έ���;�u��T��@o�ǂ�A��D-ʝ�B��X��l��X�@��p{��=�̓8$!2D����������3P��<i���Q��8є�4�=�D�A��_|��l:�Vd�� �<v'�z:���x�
,k��6d��fH�:"���	)��z���NtdTc�q�%^��+w4y~�Ԙc$���L��W�����4������b��O��'z�%���8 �x L��]ٴW�]��J�*A��%�����I�U_���fDnŨ��f��.�pˋ�����1V�c	���g��HYY1��io�PT�Q8'
�Bb�Ҳ������M&G���ҧk�"�jmѶ@�����3x�X#��9�b� ��ρXJ��6$�^˟$�N��47uΥ�Ϲ��gP]��ʡ����P�Ŝ�a�߁ ��_���1�Jz;�2���Q�S��ŷ���ߌ�.��r�:����]��d��ż��f�$�sݝ3-]t��ɷ4C:��H�w��1������a�z'�,[�F������_f%%��V���w��!G�^�җ�o{�j��[��_�g��;/n�4���4�j^/+��gN�{FL*��b���W� �_��6�c��1�S���m*^��C�$��6t5�rL��-)��{M��5�{���/`�k�]m=:L�����_��hСlBGLP���w+��C��&w�	@X��$��<r�~E��ޘ��U�����@J�dL@�
� ��VH�q��W�7�nF���5���W~�O�$�#��II������Dˤ��E���AZ8Ǩ�]����V�Sn�&7���X!Bj�VD��f@��+9(i�%f�I�$��M������,��u D"��ñ��ν=PlD�h�u%';H�6�P�wi)�����n�N�~�G��z��wY�d���k��3X�Cw���{��	��@��5�"/w�쯟l{d&�V��
{����~u0'�e�e: SD�QXLۗxkB�X����Q��;��sM���j�G�D��W�'��b��&>��u>��d�bP4���� P&���6���4��IUc��Q�����JV��ý�$)
�n�����n)�sc
NeŦE\fH�g�y�9�G���>e���&�)�],^}E��Y<�V#=�n�_�0�����۫����Ȧ 3��̴���+a�@�#N:�~�%CVIćfBhD�'
�Ô�|�n�΃���.��8����7�ߘ=%�y�qY�ݡ+��C7Y`8��ay$-ר���p\���E�\��ξ�#d��q�������`.(p+�<2��˽�V�!x���k��L��û'�@9^��`����ӽ{;N����:C�y��>,�A*����
�1e��RFPqJ�8O�5��`��$��._����-�S/q����Q<���;B�մk��31��]��� ~uLw;☮����u		U����s�0<��BX�f%�<�G������%&����>W�%T�,B�K�#���3��	�3I3�%�iO�"�`AN�b��1E�(y���=�g��ġ�9���nsTY��H?��Y��ʿpc��YWuDH��]4���i�-A�atQR��#e�-R)ɘ���.V�NՊ�飯�w�x��h����OP��Ec��{���Ԁ���-X����\�,�ݖ�# �ݞ�:�j�a�#!�>J�3�ʃ]�G֒
��a������n�ʾn�E��*���m���\�B����:ݞ7Jr�
�)}�m���<J+�b$��c[�JB����t�^ȌN�.���3���lSZ ���ҵ�~-�C�깯]�ժ��p��������p]����"tJ7N k�,�\,���7�͸����g��C��o[)nѕ�yѰ4/�Y�Io�ai5�dS��6:%i���4ʼc*��m��2;.�4� 㵛�(������k|��{�]/m.Ȁ<��mFB8C����U�	ġ|�:O�]�����̮�����x�����b{�z+���ʲj}#l.�Jl������HM�%�5�0z�ɨ����=Չ��6/���U|X*=&>P��ճ�31?X)����巼.�6pp[*M)�(-z?{&�<_,?� *���q�@?C�#�'C]��T���O1-r�ôD��o'3Z�{h��EIڵjm���%�#�������K�|��GD���!�Z���ZY�%��g\
����&c�{��}/�O�K��}��8�����')mHfns~��&�1Vޟ��:��%�����?�9e5Bz�W6»����k��зd�mk7ca!������D/��^��=,�&�
��t�����̷���y�Y�NrP�b��L��C��(���]��N9��l>��sѕ1�-,�&�Czˏ;�~U���2�?�okۢ�&���Ncܮʛ����x���
mkq���Q)��gp���-s�	����������W��cU*!�h�/�S�;���DsNc ���� �w����̘^[WVtR����w�5�2���jwJ؏+�����C[���ؿ*{�hd��/���+��J�@V����&��Mc�j^�F؂��ß��{�Ȯ(��ͽ�Ц�X{�γ4>�e��on���1^�Z{XPi�/�|�?qϩ��T����+���(�N(����'�
V�{S�d�v�_$ͻ����oq����6��fc�L;��8��T����/,�<[=>4���j�qR�����Y�ƨ�-%����d���m0&�糺]�LE���vv�l�-�ki��*c�4�s�`�1,�ԫ����� �>�ם�"7�D�W�G��]{��*��?#��}с�U�~��2-N7�Q�=/f}�<��$9�p���9//Ĩ�|�PS]X���F�G����k�9��!����@f��ֲ��!i�����������;Cz9�"�񽐲�>�ԥ���v	�,�u��2T�c|�r����U9r1�o��_J;�p���OJ��=�1��q�g�A���R0K[�칎5����1���s�-s�3Q�r�aa���~[U�dg�<|2w>U��m���8��/΋�ñm��.s.S����g��/���sé��SY���TWt�i�3gX�OV��ة����՘�6�h�|�ϭ'6�qR�)�z�#����,���+I�s�z��M�D�;�S�~�^�����|T�f�(쳷��j�x�������i�(r�YIe=���	v^�������#n$�F�sk�ƅ~{׎�7������d��[�ڄ4=��p�`ku�*e��lԋ�jmh��큮��d��:]0��MF�zi��ib�l�5���D)�Hmwm�f�Gn��B�c�{��ws���2�:\,�4����>Bǔ��W�,�B&Lw,E>��>0��9�����z��nHj�g�z?�^�$�¬S�{P�m�ELҬQ�����_������k_�S�W�<����.�3�r�����u�-+O�؞�����L��L������Com���&co���)�`�gq>R:Ye#��o��u��t �VV,� ,�I9���E��$Nn]�Z� �^A��a�l���f���$&\��D�h�"L�\ocTOTr���u���`ɕ2���<����a[QNp����
H����JxZʱ'�|�e�~�m���կ*N�A�6r�p�Z0KW�м�MUg�H1ɥ�n�~�3�c}��!=�rEq�d�d�Kki��3||�IzoPM�}H1c*sVp�i�4i�x�F?����5Ϸ2^��H���"<b��O�MH<���0��Ǽ>�z��Ы��D����3�a�q��B� U��*�iȜ�d�wb���)�Ǝ$��j#�v\_��)�n;Zg���b���}j�'����p?�� �5/ν�T���V4������݈�v_���2�����l�
��E���G��E�|�)�d���
~tr~�<���f8�p���S�j[�Q�����7�
0�B?<�Jxv�;��;��V���u���P��?�tlvƌ�[L蕖&��́�N��63[e1ۛ�� ډUʈZ�qvK�-\q�i8u�v3v+��uՄ��q��~�j��Z�)�����ZM��I���&8N��|�� �v�x=[�){�W]�#N7E�^�^oc�ԏ���w�yv��w����q�D�	D�\�#����?��{�]��k�:�-�}z�P��5�-0��@�eT#�Է��E.�C~kDy{�&�ׇt��K"3�*˨��钦�?�.�x�vD�ˤ&ʅ���f��<���/~�,E�偪k���3A�@z�5�|z�E���:@�i��t[��)1����O#\��~g.K�g0�]\0��)� ��O)��}�����
 (MD���z���7˘4��c�ffC�����#��j���P��Wm�͗�<�-q�iؿ-� Z�xB�еq��L��ڗ�\��N�c�jĩ7�\���y��Kt��E�H��'�}s��'�l��6"_�D���3�?b��i}|#8� �n;�Fr�sR���x#��Ɨ�f�#�I��F-	�e��d������UiUU������+��=YR�}����6�;o����#���e�[(�w���oݶ��
Q�j'�ouK���b�Ә~/幎��_�g�s1��b���J�p)����+*B�ġ͇��'�?�A�@ �N�(�0������a]���R��}�x����1��k���$c��Q?���i�"C�e�ʇ����.����?v�#L<[�P���,b�
 ��P�O%�[]�2N��~>��>��>�ܡv>ힲ �t�
/�H�9+��5%N�^2�3�vu��Ҹd�*�4YH��K����Z���w�ȓm{���{��Y�aa��5ٜ���7�0��R����q�2�i3�h��}�Wi>zB����ӭTV��0�$O;�ܪ�y���*Y����x���>�Tf{�a���D%-*'�[KL��Cs��ܨ~����������v�ND��͚=ɮ�o�𬁢
�*�_c�ׅ_���<PI Ç��;�9Vhjz�76�6'e�p����U�j=U�8�@��X����=>�*Z(�y0x���[�>ܹ�p4�*��`[1Ϻ��oU򄀏�wF��W_L{�"��B(5qUh�&�3�{@��5=ʕt�.��Ӄ.~���~H�
x~a���oy�7-�v�*T�G��T�^�q�-����N�>��ʩ(c����[�E�>��(��"�]�Hwwww�H��H�tw�t.�KJ�s�����?��7��9��3s-�Ar�!�5n#.�d�ɓ�6=�����kJ�2XxNH�{��c�D��dP��*x��@�ڙ���4��8����@m�PCӡ)?sQ�ʐƓgqA������������̴�Y��I	bh��+�2���y��^�9�#ܵI�_�`��@������EI�����w�}�c�'��g.N�7c؄��w���*:H���Wu�<��t�+�߀:��/uB�ٷR�����W'��Ӈ8X�?W���j�^yF�X;�����	ˍ���c�:k���Uo�v��YH/�|X �cC�~���� �74zœ?���ķ�+P��k{��l.+}�}�:3�[����!������L	�����'@Iɭ?�wW��U$}�l�=1}��	j0c��xhp�AM���Iқ�Zzs{���
Du|�="#Y�L� �Z/�����)t����g���{p��e31��D(c[�+\t� T5VLD���5z֥y;�r�k
̃J��
��~��cT�n���s�&Q��F!��"���C�j�@B�L��9_,�h�T|ꌻ���a�N��f�j���W��jiB^�������P4�8�8w>��L�m�W������8�f��Vԁ�t�G~�ກl�����G��7Ѓd�X�G?SK���	��ҶtO28t���Ԋ�Ȏ���½��������FUh�:�=�����ıi���Lh��-lI�+TJ�(���#�C?��bY�z���MnU��)��a�d�}Ldn��z�d�����g�+;�C���9��kJ����\@�y^��c�oX�#��%����Jet��u�M��rk~�d�jXG�*W�Z���Y�����"!s 5�G�!��
`_��"��q����?>�I�H����{�����)(��=�OY�+��Dy�;N�������`�,��2��rS՚U����)6{<�M`��ߩ����v�o���zkG��'u�H�������Vf@�E*�Ǭ�F���B��s�d���ij�[�ּ�Z�c�M���c%�Q�]���ۤ���sܟ�������)Ъ�� t�X	�9�f�i�z��φ�|���{|�w��籱��K_i����zg�֩˃���ƚ�r_c�K�[�f��r6�
�ausm�d�Z�^���=-^��D����V]n�����"Ni����6-��dB�Uf�����O�,C%�Z�a%�� ��� �����*��څ�|�61k����eE�5v�e���q9���Q���/�xG���ݗ����q.�J����UPO���ԯ�?����&d�<�	�Lc~\�3��T����hr{�0^�'��A��~��B�-/��K��2(K
~�ɋ�d� ��Z�CX�wcƖW0�3tT+�!X�L9j�!��>N}5VD�R���Z]	~�?��$�#f��U��n��
�l�j��4T,���F��4� llWs�U���j�O��ID�7Zpfr⻚z��4@eS}({@{%�^�ymt�(`}4���:���H͌������\��n(�8w��@4���	�=W4f���'�TaȦoC{j�<ҧ�W^w/���BB1��аq���Yj���sFB�Ԇ����F+1R�8���������`� r*�ŝS�1R�?a�Cajн*I����4�j+������Cp��D*M�c	�vTl��{v�����񩎟��w�[���Ų�'�pz
����l�!���������m9��Y��q;;\���e^U���E�22�V���~��Û��'r�a#9/�)�;3�Y-$� ��d��Y]74��ΪTTg�-̶�<-/�<0�78@�R*A#_��e�\t�[1tF��}�+�C���&p*���8����JKN���(��plͷ6����}��ڕ9�i���;N�� �5��VS| z+��Va/��+'��[M���[<��I=���ߥx�x=�l}�X�C��;Y��5V@-�JD��<0A���"��Z�=���.��g/|�"��3��r�7�ѷk�� z�H�XUnpU~�'���+��ɔ+k�n��C�I�Ö����.�q'������kw�����U� kk�q}���tҀٜ�/ᡝD�R���d
�
�!�C�%�4��SdF&�o���.C�ߍ���rO�u�0t���3e���JQ�q���f@�*�t���
��������P��}�v����E������R���Z@x��zm���ek:���fʏ.�����d/�f��{�Y�ur�h�7	�!�|�V�&�� �tB���i�rq2͊E�*2��0VEZ,˓��9x���\C�dЏ)���<��w]V�(�yNo�gp�n�s�k��n�n�}��#�e�-����W��8�@\�3R
1��h�oe��g�kA�)�p��H�t��Qs㆑==_p��Q������)ee�p{�^0ۆn��I�a��U��$N��O8��	wa�-È���_��V�[�)����Xܑ|j��N� ��}q��L��t�@�����4Z��8��Bm/�њ�<���,`�V��#��������M��5_hXfO�.���[a���M
��
��W�@6J���Y_� ��n8P&]��y7��"���%�m�������U��]�0Z	BJ[`'��G�:�	9e���I�a��ڌ�8���c�I�3;����״�m��*t��~�>�|E��W����r_��q&q5N{H��ю9~����4�G��?S7��?��BvIQA��σ��ݽ=P>��@n�'֯�����͟
�5����Q�W��ƫsN"s rJ��;dG\�ї�*A<���	ruQ�r�WJ���.E�	�=����4G���)�#ψ�=�t@��Ҝ}�`���r{*�*ù����{�ѵj���h@s�����ٷ��q*�݃�4d�״�����W*��
\q2���ί �����k*Ö0���
���W	Ԭ�h.n��T��Cb��}�(���5'E3��$��?����M�0[������uzAKh�?*�3*��݃t���4���k#��q�qA��vf�;"�o�/�"�Q�	hx���V�$RJ��T	���F�u�ӌ%��| ��J�!�Q
W����t��Jv��ȍt�������2�3g��������G�c�l���ex�����W���p����f,�kݥ#����PO�&�!)7�Q8U�2r��C%�շ����R0�.q���j���G�����Ucr������N�谢66$' �қ]�,O�z�w��u��·y�>����s|u�^�H��a#DQ�sU�e�To]rUO�YТ�����H����tt�����Q'�!{�6A'����A*3ĉƬ�i�C=39��������)4�G��ǻ+[�	�u@ n�2N���8(�p�](���˯yt�e�M3S��Պ�/w6;� ���6%\}�w_�4�mٺ�W�P�fV��'��y ~y0Ewa���=R�q�gW7z������ae��c"ѫw���h�?ƥ�Ϧ��.U� IT#NYh�ɣ--`�������W�:	��(~�E���� �W|"[Z|=X�&]7� �x ue�?��p�H9��e 5p�@ha�)�����\9ΐ��HJ�,힉�B�MsAxyN�϶qw�:��|��p����\pk�
���Fe�ۤo(�	�S �Ɲ�Na1Ki����o�Y�|29�/�kG�W8��|��wq�V���~�����;�K"έ��M[n�:�*�~�aoX��Z����{U$)���1��<E����\�2{qO��Ǚ�&���E�����M����I裯��0 6TH�u�T���00Y>&-���.�P�5��q���R�_�!�i��8��X�$�I�	x:��mDң'0:":��_{�]�`�\�En����Z8j�ۧ&����3���ۀIbc�Վ(O 4$^qi� \B_�E9тk�%�|��S#2����)˳i��d����%<�v�RҖ��it=�NX�D6��<�@t�/NU���at9.$�;�.�pk:�I}c�byV��;K-���k�d:�������~F���cK���@�GȖ�u�����hAJ륿��l���b�}4B�(p2�\��I$O��>�>�b�7
�w7}�o��������1)�D Va4,�@X���Ds��^e(~���l�Z�WMD��� f�]>5��l�hx� 2�`N֩N���?4�خ��I>�Ur�����~�@W�/D�M�t�_���<̶c�ڶ�� i7�U�a�~R�;�u�+O���I���/Z{E��] ��
���1jaL��S�M�&I���g����s�w��C�{����y%x�AΪ<����s��2vp~��4���`��U�;��t���㑷��R	�W��>��g���Q��P��׆t�1���<�ኍ���$#��_�zFx\���T�nZ�3��5̛~d�ʐF�Q!��x�]f���o�����#a!n�2J\G�yy�]�~�&��'�m�%�7��� �P�E�����[𸨈���`xn�����T�_4��q�׍<Mʖ:�7,�ˮ���b���pұ7~�ģ�={��S ����w�l۾��懖���7~��QQ��u�u��@��*e�IK*���Y=�x��꧖��kD[:[�C�K�Z]TX�����@G ��)��X��<Z�&&�x�݀��؏3�3/��r��������E�(7@g|��6�(lrZ�W�@��F W�:R)�!���S�hL^R�/�ѳ2\�=�K1
�Af��dL���DĈL���_�ﮩf�	 �1wS;�N�2��_mQkO;	cwFg:��kܙ�پ��5qZ^o>	�o_��9�K����udT�#	KP���K�ihy	�Zi���Z��������;qF#䨖�~��d��@DA����hd��u��������A�P{�SV"�yl�>��V�1@���k?@���e�q�+C�:Z�Q�S�E ǻ� �vxs� ���x
�	-��l�GʤM}!���F�q��'6���4�����~��)�qql��Vx�OTx\�A��_�J��pS���=3��;N�Z���dZ��Ądh�Z�� ����!��N���J�D�/����<���ܸL�=��#��~i'۰���h)�j�o���p�N<��"���>3�If-���k��g`�O�aq�w�HG�-I�>31KDB��n��@�XE	��o�%�����}-�Wʭ�S�Gvo��`.5�v�o5��|�}jt����N�3�!�ip�nD*� �$n���hn��I���߂��,T��_c����B��Y��� z�b�0>�o䌵v��M�ew8n����Jc+]�����>gG���Qڗ-��p9�Z�&�Ą6�T{�����dC+i���+�]���39ύc�Yy���1�Z�J���^�����ܐ�~|.������wAZ�ҳ�ͫ[��h�/���[4���d�s� �/�/�l~l0���
���T�k+�"�DI�!�����ھ�^�`U��0K]d������e`I�̼�8W�Avi`xOd������^ű�D~c��`��\HV���o�vu8�n���j��X)�y.�JI?x�S� lo��'��,ז&P/��A|m4��u�	�\���T�K��.�:36�B�в��K�v��꺪pW'���Ru��5M�Ζ��c���TtEeVn�O����%�!̛��Ld�	x+9c��R@8D䜨ن�7���/�e�\-8u��<���#ι��q�$x�;|��ydޙ��'�"�2I���6ԫ�Y����EF��5�:X|�ݣd��V%������]�E��a:�R�V�����RUO&Ĥ{�I�Y}�j�K���:��&x��������)ĵ��@ح����ؗ��}Ȅ��U�++����/'���a'�4�d�\��w?ј���~<6Dܱ7�.+��'�]<qAB��3��+5Ԝ�W��< /_�<`���\�Ӈ�!#����򃓍��H�|�}�k�/WeH=�"n�7�6�;W���WL�5	���E�"�N���1�O��h'Q����S� ���AU��BT��+x�ċ�p�o_�3X
O����[
���4�ߐ� �pݸN�N"睎7I�#Fo�y��BA!����O�`�����)������P@�b�s6 f�KqB=ɕ�:D��ē�v��Z��+�ү���F�z�&ݿ�'�y�̃�ٚ���	+´P�D�lv� =ǯ���OR}+3m�V�2V"�_�q�o-f����*���l�dv�X����3��������Y�RWtCP_!��7@���dnٶ��L���5V
r�Z�F}K�7�.*��.���O�Hባ>@I�����	o�E�K#)q�5��ك��n�ůꚨ�$
0�]?���䚖x#�c����6� �<�m�#�/�C�_�Ju�MhE;�;=2{�/�]PR�"< i\�j�wɲ���>�(\�����g	��<��k�p������h*?n0l�\C�6g���w@et��h\^MXD8�م�d�v�k��ۼӹ�֥zgn���+;t��"��q����V�6d\�4�`gtɸs�=����&� ��l��Ҽ��ZpTa�Z��n�A ���ť���W{|�?	�$_W�P�xº�d��p��xo2���cSS_.X��^��g�E�J0\��C�C�_7�osv��s�p�uWrn,O�H	�w�8�T��s����T2�u�*��[z,��v5���}4㞖S�>b;i��^��Z�w_�9��f�����M�{��>9����(8/Ǽ��^G�/I�(�����'єU�7��ʖ4��>��5�?� v-4#���{�Ŭ��]�"�{ :>޸�r��Q4��/�F����̎c�.Zky���XA��[mG�6S�x5�q.C�Kz��W\�t�����[�"�lXף�i��&�_��-'+hM Td~�,e�q�$��{$<��𛺨�>���}`\3x�k���E��}4	��b��叀���^ovd���OL��tӈ��?�$�.B��mP7 �ۭ���ix�VϾ��%�z������^;n�DM�05�}�Hh���	��kG�+O��-���V�!ϖљ��6d��GJi7��u0���"�Ս\)��y���{?Y�e�˷q���4��
NGjv{��t9�p�+�ScFj$Q��Km����{ �I`f��)&F��mӼ��	��|J<���M�mSڕR�@���W�x�n?Զ_�*FJ�xd�~�d1#`�M���+A\�1��Ź�;�5���r�%�S*�'� ��be��%�]��n熆�� ��B"��ᓲ6b���
w<� �i����[$��ߥ���＊KP��I�0Kq��&��?[<�k��}F�}
_�F$�\@Єg廌��vw(T7�	Q�-�ﾭ|�#+w�k	>���e�_�y]jTJ.��[����_�E���CX�?����pC�iJW��.�Pw��i0H���trRT¿;<�-��Ys�vq_կ�K{q@W������L�C�PE����7淋? ���@^�A])A�|ti()(F��9����,[=ܕJ��|���h�r�0���|)
?�v�s���� �@W���}��z�_j�D+�,QĪ����S��%�!��ׄ_ׇ��u��9�m���T\=D��A��P�
tQxG�ԝ����P5�*P�(�1<��o 6)�-$()��j�4�?UVRQ+6�;�#����b��bkdp(��y5#�	�k�u�pn]g
��ŵ��X��U��{{퀿�`J�ʼ���kH� E�߳&���ސ���ȔwXkCCO���bj�x�]H+�~���_v3T����=��95v%��1��U��0 ��O�Ap�t�D~��k����u��=�: ����qf�f�B��:�f�7��F�༏�	$�Щ
Yu�b??a����2�A�f �鋁����J��ͫ"�2��˽�|ߡ��������kÎ ��3�&����ս�����x�u<�v�x�\��[��N�(��]&b��ӵ��m�[�k[�9���2싛���d�թ h�_�BD���G@�)<�>�=�*_��N)%�/�h�4÷f������"�]ģ.��%�?q�p�Eg�%�|�Ħ�8����@�=��6I�;�E?� ���+�����4�T@-�f��2�`���u�o�(���ֲ���<x����{Nֶ�1^�UESj�p���̬�}�� (l��������I:o*F�yj ��NB�A���#�B��Ʉ��%���h�6�G� �$��dq�w S�Ņ<��(h��@�͢}���B=8�����aVv�/�]���E���.^���g�gq�K��ۀ3����=����4%�g���lG{��� h���m�pd׸\FK��9�(C�f�Y.��"�`u��Ʊ Iȴک��ȑ�實�<:ꊅSE���lH.�w@쪍��6�@��T��-M��$���2W�e�G4��SX��<B���6{DWޯ����a^�-]l�Sh�*n��S�
~{�_� �U1�x�������� �(������>�h�qC�����ɺ9���+��U��Bx�~|G�q�p9�O,~>oYe1c��gYcf�x���Prbrr	�ч��Z'�#�@r::�N��%8����	c.q{m�O��VrJ���
�D��$g-�Ӎ����A@���L�������DV�0����?�7�pߗN��p~X���3P
~���M���B[T7������N �F���>g]��u/�& �A�̟`+K^��@�e|�����f�ij�{3���jb42���`CK$�Ü�����M�7wx����Ņ	�ײm��]�x_hIa��c����A�r��X]яߪ� ��+�������L����a�ڇ����B�q_ee��D��/8�����G��%�η��<op2D_�������Vd}��mf�:�X$*Q�������[i\k]E�-��\����Є��_ND�Y�xm ��R���+b��9���\h�U�+��p���}��Ӕ	��6� B>��Jz	��K~�t�'X��L����,��b���_4#�:��&�+n�VyZ���NW���آ�ԋ��=�TV��[$�GO�3��?H��ᮊ�����]�~����|��wuJ�l��ٳ4��� �PD�$Ȁ��]Q�N�:��.�F��mp�6�ƪ��H��*��nq2ј����Â[��bJ��Wn[(�0y��#m��	�_ߨ����C���]M��m2��.�4U� �Jgܟ����k�7Þ���A�m��m�ݑ���g��.(`y���؎6H	�D������b��|xa)Tak$��)���rXއY�������:(�@W�ڸ���h����5���m"C������9�[�_����G=���.͠dZ��Ij%������a����K�A�}�f������@��C���Y-��'z"p�+��T��sՖ��B�w�c�!o����zoE���!?��}�V��v,����&:�dṍT��W�0����}�_�87���#k���s�4�عa�M���]7E]�஍bb�UC8 �3w�� �8&��ą>A��.m&Mz�O��=&��=w�����*T	H�ޭ&F-g�Ç�cT��:y�
�/��J�Ĵ'����j��4�M��݋���hJ�رL�ɠ�Ez�?�mr� �&��RѵY-L����`��r���ʛ��ӻև\�c#�DI��o/�*� Q%<N�(�^c�������D��uY	y�A�S�����u�mȫ��ݹv� ;���8��^�9u�'��?�03�,�����У��8H���3u�kjsڭ�@�Y�vM� �t�vt���9u~�	�
��"��Q����Qj�ɾF��y	�$�_h��6����x���^��'�e�̡k�y���xh_9s�k���޳Oc���W��K҉ ���Q9�� ����	ڝh���Y^�[�s!���+�(��wg�cϿ�T���͆^���h2�v��1
&�mw8��[:�J�O[����"@8��k��>+[��2n�,�/�Ճq��#�&S@�h�<+)+;HA5N�_ru��+�9�&Aü��-Q@���t����H{����� ]T�o�w~�&9�n9���tU����.��m���FQ
�m˼*莯�J;i�Ze(Y @�����+cW]<ksNΌ�g^P���j2UPi�.^�"L���k�*��vps�~CC�[W��_�y�7�2��AJ1fr�/���a�~�3(�Tpm��̬��t����A��S6��|e�=S&Q��XG�.� ��՗+���>���̣�m\�p�ձGҸ`�'���7�9�g����X @ 4jo��_�g33��nD_iWKf �d����ϔՊLxul���ֳ�'�|�G+���̔Έ~\�����N�3�X1�@C��\8�3<\�8�1�/{�I�5tK��{|s�x���ţ�z`I�2O,Ȃ��� W�ɘ�kn�B�U��Դ�����r!�W��>Z��q����G�O�������$*?V���M�ղ2X0]K�s�OL"h"�`"R��g�	>��N14s&{jS)o�dŸ_!b��n%Z���J^u=��msx�}�0��⾒�]�k A2<����k�o�5�CҸ3��%>�ۉ���hP�=L�Q=)\�M`���s> n����5�����"��.�,�����(	� )$	M#��tȆ�e��ӡ�`���<�_�:�N�+*��Y�){@s�`�^>����=�'!
�<��*��Z��竸/��������hў�^_x]�6rJ),jj��y���i�����ک�}��N�N���w@ů�X��A|�-ߥ� >Y;O����e��\{0%٣]�E+3�>���n�xP���Av����Z{Dr��F�Ʌ��)Ǜ,���L��gT���2~_�r��݋��j�<����<5�Snf�Ӥi(�Ŭ�5f]\kp-��͇��'o''�;=�I 9�D4A������e�������A(Ɇ�'.m����_��ݤ��ܩ�5)Ǣ�)i�,�F��Wk��#)A�m����u����XM�K�l�!�[X[[�x��ƕ���q�iÙkYܟ��[U�)�A���H� �N^6);2!@.�:��2W��2����]��=FP���n�pk�W�Bgw�!k�A��I6NO��B��t�%T�������q�ۼ�z9����p:�K2<i���W��}����r9d|3��?P�������}����B�'�!����L���tW2ˉ�YIe�	|�1��{4��ք������`�t�/P�~j'�YCl�6_͙��>�512}z��`2����\�9/��:�����e�p5��n�;���L��ji��-d���!x��o:�OV��̡M
ɴ�����B� U-�?+l����M��L��u��z�g��=�z6p }x��p�)�������R.�𱱶�9�U����A�U���I_I_�AԺ$Z�r�h��|ŦǾ5�\ݒa_nH��n�q���Ж��/�����k�oa.�'��]��,dz�oddyV����/Q"� 3���~��h����� ��p��y�E�b>�L�ӡ6ͻ\��Q10~�S��n4x���"s-� ��-+dgT-��}�|�a�����h ̗�~>��b!�V��eÕ�3��A�/��)O�G7>�y���g�!�g]ܝ��|��P&���;�R�T�v�,��Z���m��C˳ʋQ��	��&\������ֶ�n.��[%B[�&�/dW�?���P �G�/ЎQC	+M�Z�����<�eKkHq+`�;|��U���T�[�|�0�cò?*���lS�}�Y/���l��y���2 o���z3�rk0��-��V;��I���R�L��7y����ב5��/Jx����pV��9��@��Zھ ���۱R����>�ߪ"��sg�P��i��t&R��~�tɧl�R5��w߆.#������	���s�;)F��D
lN�殼5ҕJ ȧ~�P����{�������5m��r��i|#(���:��	� ,I��l�_�H����o��N�U�(� 0���jz�mk1��"wكi�gF����$���&\'��ۦ��()Y�_ںI�_&��YK�=��CJ!n��l��H���K��xG�������t�&D�!�y���w#�HN{!�|�ʊ�8�����Nky��شj��V�*��=p���^���W��V����~��*Ez~y��%Yk"�/�q�:  6�$��(o�����hw��G����xe�)���o�mG�|6q p�	M�w�?�tw�=��W]���c�*�2�F3J�g�D�2�w�Ob���}���G�ܞ��Z}Z� ����~��~��y���-�U֦q4�϶�ش��-L���@G	�xQ�K��%MgC5�Yk�+����� XhFk�^O7Ϳmy���$�F�2�Y��iЋ��zni��lu���@a�iD�W�����ډ �[��	��o���2�H��ѓq��'�Z�$�"�	٪׹s��Ӟ�T�06"��p�.�DA�I�-����挏���Ť���K�BT���K��!��<�O�4W�+����I�6l/�?���qc���C��	2��(b=y f*�q��@���͖iZ��4���q���S�]�cg�H�K)<es����F؁\�^'�Y.`�EG�)��Ĺ	�w��笿At����V2�}�}��li#��kITT���ӥY}*TS␢��*�D2�x��@d��t2K�����z��aQ��s��{r-��_D,�l��	�y�$C/V&K[�}ݡp�����XW�a����g-�җX��L�]�����?	�Z��ҠJB^d؞ˋ��M"�f���EWc��fae��2����S2���Μ���A��_��'곡��z��C@g�#+<�rf����Q �
Ly��1˝�D��P�ڸ��k�6a��e3�S�C)�Y������?E�W���]{�8u%�~a݋7��,:�\����0VQl;�c��ڗ�B)�=�n|@#N�kƢ�=?6�0y�v�c+�]nUfo ��)�z�,��bhl͟%<J�
�\ i��]un�Pb �"p���B���MZI̱w�@���4�u�Vku�.
)��+���s)&fod�r����(�n�z�lvЊ�����zf�0^����ԏ�O�a�}�V�TE��f�t%�ǈ�Ih�%ھîR~�� ,��4���)u����^[��A��ssW�����~ɜ>����!'��ßta*�]G�V�F6��)V?#d⥈ȡF�T���u����������?�3_|�J��S������'u+]�9����y��ɿ|׭�ݖ��:�?��!���X�D�%nߧ�铇·:_��vVP���H 1g]*
�$pV�g=��1ڟ[�Ę�R�sB.B�w]p$}��G��v?�K��NҴ���L��{�	���wi����ۿ��sD�D�7��?z���0���D�pcK�iЩ���ʻ`�؉�~�׎ʁ��م������a+�[?W�V�Iw��Gp���N��0��쪟�Tz�Y�X��������'��8�z
:S��L�	����ьI�S&$]��&�CK�W��$�Yy��������p]r㥴��
�``�Ud��zt�yo����Ɔ���R���vi7�!R�t�Q�	�ҬiQ4;)����-}i�i��e�gc�I����	^��h��8i��U&�jȕ�|}�5ZQ����K(��\C�t�i��پ��}F����F�+�qL��H�F1��_���,�L�]��c�E/�����,��8�(��4d%��C
k�\���`���f��49b�.M&�O�倩d-ا��D�w�yC�&}Z׍u��Y���c��̃�q����6Z%���#l]�u�ꜫ���s���$�9_����k��S帑&ޱ�2�� �N�ҧ�4��G�o~��|�L���["=�j�y�Q݂W..��u�T�P��#�k�B��Gw�Y���'8]y�~����0�W/�h���+P�mN�q��ע{�KW�t`������?���f{��ls�-��
&״�7����f�0��ܢ��IS((Z���s�iQYH1:���Q��1��|�3PG��Q��Z��/�O�)�YF��i�A2p�D�'{����t�����Y��v���*���J�u�zj�&HXb/��!��{��iGd���m�%�'Ō�B�i��h�5��0�0��ҭP�\+^��lVh�\��9�0�d$��ߨ��.�$��w���b�C���/F��t��2|B�%Ĵ�#�/�����mwwd��P�@X�0�S�l�ĝ	�4��%�d��۪:�i��ڔ���k�nSFB���2�sr"#��Ø��H�s���{��F��[���e���~ʿC���[z�˒��Pb�q��c��x�����S�ï�:�^W���'
�q�J��ҩx�g��'��f_�,$*�a�ZQ�����n��L�"N���>�uE䞴?x�Ǣ�&��ڈ8>�2\}�s.{Ü� ߀�`�w���ݰ�����9����T�Q��v[4���*ؤW�2� �`��}'~	����>5�ꭿԅ|���s�E��s׽��d���N�c�#G ������m��q�-ЫX��AG\���/_�!6��2C�?��sS|���ygJA�y�m��+�G\zګ��S�<���\Et�?��ފ'1�M�����XOI�g�d]X����˒��it�Ao�~G�'�·���jg��[����-No.n�<�C�&�]�~$�g��=���$yo�4�L$_p�ϝ׫��^L*�Ol~F���7�����s]�^�,��z�v@�:�>�۲�>��R�f4d�L���An6���w�Bk�K3Vߙ�2����y��G�ĭ� s���Y�Æ�c�Ŧ��0����;6̚����G�|<3J@$r�n�
mT�ދ�}�z	|z�?���(�=��a ����2T��C�l~�Ȉ>2������.S.]�2���\�����>��n���D��a�����L�����%�R��w6t@�����M���G}g��WO�~���P�>�b/@�֬pW�P�%nT��w,��m��ſ-��~���L�q!:�j�u ��tv�����?���߮�I]�q��񦃞.Я㒾���r}㽑��dЮ~�Lx`3m������7Y|,L��6j4��x^'([��F�\�a?(�<�oTwf��*���	��F��o6��ɮ�]�n�e���z�B��/��t��������־���ˀȯe[��l@�v>��,R�������D��bgl]??�Z����tm�Fp�\=?�>?�z��󪞸byEH�&�#�c��0eΝ�8����� #t#á�;W��Ŗۊ�#i ����3//���)ym�7�L1G�f��Fy�o�7�b�sx��	1d�]�3����Z	���c�$ٝ��X�a¿`*�I��q�T5d�:54~r1�p��]ɢWb����V�N��"$�t�p}�=ީZZ�Bh�'t} .��D��ж$b=�)y/0�L�i�[�*�u��ֈ�"Tӽ��b��ZN�1���XNb�aa>)@\XC�3���6�lPY'|[o���B��6��ȁ���wR��}(�/7o�[yDݾ��
�:�/"�'�3�-|^��`�"H�b(0�|��95�
�#�¢�ަ�L�[₧oHO+ޭs=�ENAh����.������j]�"#ꐙ��sv�lG)ԘU��"�鏜��&���A�o��<Z���^���x���+�(�2��O��z��Jȁ"��M�2�gO���
����� �L�tF����h�0�)$������l���0*����.�?�*�ѓޯ�������v��&f����w��f�S�>�0�Z�-�GT�Q#쇟x�{�9%G;p::iV�  Ym�^<�W��jǒ ��o0������.d�h���Q(F����ڐ���a�̵�x�d��R��G� �K�RS2�oj�=()�h߷|�#z~/����T(�NSuW����XFm~a.]a?�w��L�{��˖� ��F���/�9�f4��GoIA�oګ��w���X YtZ���u~B]��:��"J3lp�b�vƯr�G0�Zu�5�����T\n��2x���Ωh/�^��Ic{�'p I@U�F��t����]m���$�iŶ��
0&���k4��P����e��al�$x��w��m��L�4ô�kd�ޣ�����Nf�Zmk̸({.\�YZ�<��p~SN�\^��gc�ɹxF����Ǆq��3X���%zU��j{��g6�/�_�;`O��m���BKj�Wp����빤���A��d{����>�'���VE��9S>{�r������@�� ����5��ӵf#ٻ<�"��cQ��;ceD>#L	���3�L�� ��?�Xp�>��"4�� �%R�5�0(`�ak�G�q���i5�+9[S,U6b{��B�,OC�ǅ%�h�l�^zK�χ��r�Eg���>L}��~Z���(��1��B2�E��V6� �o�@�����.��@�V,ph��3�N�\w	������m�Y���x���vh�놥6�-#��Z�TA���"?��:�h�����>e%V�t���Ȥ ̽�$���ʄ�G؀��������F��������K��EZ@J$��n�.�����A߷�Z��#k�y����o��_'M��r$��!�)�M\缜�Z.v���j?�]��NH	+��Tܬ��T&�gH|�Y�;�(;�n�)Y�ޢ��tU��+��Ҿ�|lUH���H&1Δ���hX&Oo4^�Lq��P>^��<qx'!�NqN�燬����F���.ý� �[\�&d}�����R���B��Qɠ�M0V�}���ؖ{���(5��0�b��|3������ʌ�j�J�\�p�,�wz���H�+g�t���W��e�mY��N<���W���:֥�Y�ur�b��|O��8rR��GM&�4��z��lǃ+�h��ϝ���=b�ֈ�����FETiQ�&����\�Ye�Oߥ��o0�7��^�S)AO2��œT"Wp�G�& eZA�>��Ppmk�pXl���Ge��|�f�$����w�ܺ�����oa5*;�*��ta��� ���a�a��E�u�h�d��4=js�5��0}-_����>޳�J|;�#'i�t�sOa��b@�:���%�d�����W��)A���fy�~�g��|�y���>k���k*>��'�a�e���E)��wҠ�� ���'Hh��Bt �-,�}�2hW�j6W]�p���>@3�����9>���t����j<�^�X�"�+"��� �8d��S̎��ږ�|��\"�Aw�n�mO���z�����6ԍ��ʆUK�X��������Y�<IiJS:��WL����l���-='���b�
Dr�J�u��{�޽����P��\[��������n�����S�Zud���)*}�ŵk̛:�1�^߈��*����o%/�m��p�s]�R�Q�a�o/Ps�_y�Q8��Cv��qm����U���<�ˬ!�dQ�8r"}��^���E`k���9\�����>Q�X��tԌ�|��4u ���[ܶ W�E��QJ�\Ũ��<e�!%0|E��Oq�&�w�DC�ۮz,j��7�D����7�x����~�����x�!ZMHL��|��SA���8:�����8n6���ک��V
����2y��������h�!����&��'m�����;:�-:R�yέ8L \��I�u�e�d���N��.B'�?���,O�?��	1�zc�8��(�?#G@x>���[�5����\du+0�DW�B�l��wL:
;�m˸A������+�h5	p�@��
!^B�15[���[�t�Ł�J����&/B��V����&U _r\���☈���QƀZgg�_
��o@ſ.t��}�#�2�g����H��;� ?1oY/���P��ޓ������`��*�C�)��r�͑w��eFbϑ+�I��p�f���@���S^J�H"��I��or�{\B>+���I��Ms�su<n�]*����
�����F�tɻC�_����?�'�%�G���AK���ʲ\:C�<n݅�v�לɢ�?�Ԙ���s���ۂ��-��r�̞�o��ٻ���q�6��=�O������3z/^���zN^��p��Z�,���Ҍ���Y�RT���<1����Nr��%ҝX�`�"}���M���}-:F�=%Y�[�vʦ�Z�:��V�����?���`ؽ�=	����]u󦮳4��o��Β=F��֞@���K�I����S#������^
(D��������t��%�+	�'���һ�т:���J{��H���̯\WK`��!B����DX9 R��d����������$m���nD����+�m�}�t�y$#���f眽D3��&��ҷ�z����bi1��m��&����.�d��^�����W�1t�Q2)�A����\��"����"i%bx�ۓ�-�,����(p��&�H�ֺn��n)S4#f	�;��U�CJ�F��P�	��B�%,��i��s�����!xԧKǈ}ۃ_�_}���5�^��K (5�!��<��K08�y�iҽ�����Me�h�9�7+�d0j�o	�"t�'����=6!�^�T�o�2���~g�����O����Pb�|�P�8{�C��W�uнk��hz����O�e��Vp% �]��:�=����O�J]���k�H�j�Y��oby�кf�޲��P�n�)��L]˦�Z���CF8m���t�CӢ;w���V@$�~b��I:��w-�B3�����C���i�a7�u�A+��Z4��Q�H�ToE��k�r���vH.J�t��Û��l1��,X6ʢ&
ۆ��ߏ'��R��b>��!�[E��q�d�<lϩ�eܻ�,7[r���dWG�0iI�\�ދ���5�DP ��o`%�vx������x1}Ɵ�%��
�4<�-��C�CAR����`l���ã�{�jyH��+r(v-b@������_��8bY���̻6��-�+ bm���?m.͠�g[��+�1a������<�)�ߎ�.<�%��	����Z�I�������3Ǳ�!�	/�P$/<���:�%&a�_�6U)�!B+g�9^�r5�wZ]��ճ!�l[���ٹ��/�}��3�0.w.+z��'fcuRz�ߣ�5��LUlϚ��U\��*��P8�Z-�]�4���G�o�]����V$J[SO�����zC�U/t�j<~��l�[LkϏ��d���a�,wj��L�Ȍ�%�E�)�W ��M�/R��%Q/
���wG���k�����N�#/G��iN��8(�@fR�"��S�w��/d������V�#�
�)BϨ�r��W]:�+nT�~K"c�Qm��r�E꙾Iw3��\:Ph�¸Kyr>��$"���~���*�FĹL(����~�$����\��ĝ$wPw���FuO������:Mvj�挕0=d�'���e�GhH��ԵDY�_%_����j���/c���%��eo=��L#"E��j��-V�g�b��_K��3��%N�����P��t��Ɖ���Rٖ�j�O*An��0�Wh�f�Fs���ڵ�}�\���r�n`�%�c"��ӰāR�������������?�{/�nxA�L'�&Ô��i-�8�� ǍC[�t;z�9ƍT�(q5��W��޿���<��.ˋ��iA{T�rM `��qnؕ�0嗡���l Y��Jq ���@���+$�ɂ�V����1��s��c|��В(ϰ]'Vp�L������|��ݛ�)o���Ս���Q�n(�y����/��ŏ��L����7�,S.}ޭ�L�z��d�m�/��>'�k��^tپ�N�$�m�ۦ�mc�ӫi�\)T/�<o�\|�FL3�{%>��W`�y�<���T���-�A_�L���z�B�]L�n�?���E�%`��w��\;�a0�l�z���Y������9��ɷ#�v�����P�Iy#R�W~RI��p�^[���9r) Q=�G�><d�=�l���E3���گ2=r~L�fg��V��<BP�B�x�F�匠0��`�*+�/�)g�iC����R�a�[A�fU�j~��E���"�� ]��F󓕫���у��vr�*N���x!�^�0���[:�b��VIvtԐ�S�x�f���3uL�S!�*���ɰ��l����[��~�/�.���2�������<�Q�0=/�\ؗ�|#�M�'�W�S���	P'�m�6���!Q��j��(�	����Kk�N�0C�|�o�
fTtK�ԡ�_���-��ڜ_6�|F��dm^�q��Ujh�,t�h.{4�s�}Կ����9����XE���j�0ckϳ�,�|���3{æ}�P�t˦���R��ZZߠV�5'Gg�T�۞��9O
nS��,�J�s
�>k��}u����9�|���:Cs�|�W���t�n#�^�����M�X&�Y�����Fn��R��A� ��,�1�ާa{���pJ ^���Kk��F��� ���toM	|~�1~�Q��-��Ȱ���x�+Ջ['���\z��sq�����E�\٪������k�sM���h�4K�����S�BIh�+��O�cCv�e2CS���42uĜ?a��$��+�$�m�h�B�z��g6������K�XWQq�^sȅsB��|s��6��fi�^f��52k���'��UT����rsj:w������=btlҐi��Q��=�G�����"*D�q���e�K���KbZY�t�r5���%dRtXԮv�s��Ç:T���CR�Ԯ��������3@�J}���`/ۜ���@^��H'Jq�Hiw���$(��ai:����Y~��v>3����5�⾰�(���������B}��X�tVq��̅*SM��I�]M� f���f���Ք1a�Տ^&欞��Y��1��qz��e�S=���ao`�-⿝�!����T9W���E�܇����/*���Go`/���B��5Db�+ep�J�|�k�]0��{�[CJ�Z�A��T㚭�?�^6e�1:�O��9BH�0^SY��k,����~����V��n�������A���m�����r����`�f�Xߪ�z�o/���6���"D�H�[o�|4��s�V����Z<��ꉳ��z��PV/�9��J�TG��޲�O�X��an��~�l��[� u��W1A>�`W�/����H��|=�t�q��Ԥ��l�"FG����V�"��������q�}�{z�-�t��#챤�W�|_����l�s���T+0
�`].y�����6�NͶ�;+d�<�6�y�)����M�����-o94���r`=潜:�==����\���C#�)C��Ǜ�U�F�-FS����°W3�|b�<�
��fbh�̥�^>�z��v� �Xq����yO*�p�_XKm��߹�(1���Ɗ�ׇ��ґ���)^�A��>�Xx^8I	�@H�>y=/�x>H��z��ޱ�v۪4�(�Wz�ٔ�>��(�Z_؍mL�Ҝ[>} ��=&�ށ|/?}����=�{`/�i5����M���N&���gظ�*�a��j�h�zę4_�vf��d�ƃh`5��KΨ�^��'���dy���rO��P�Ì�❑>�=z���'�za������z��� �4�b5	��ͪ�{QF�{�*��/�D�6��̙�\T���p�g�}8.,����Y�1�/�^�2اX��/9R*Uxʤv]kW%��~$�}���[�/}W7����;��*��>	�+����'T|@��T��������|U���&�M;X�+��6��{� j(�w58��R��(ַ��؇��1����WfL>,ߑU����ﺜhS*����ei�r�9����=|�S`^	�e���,Ӑ@>�+辌����RR���͈"�[b���הH������Z��xfr� ���G�`�y��V��T;��+�i�X�J2����<�����5��k_�?;z��.�u���� �ø1�^��߃�����3��߽�YE�('W�����@����_9k�iqdڈR���$E�ĴAC}�*����ui��j��j��V�L+����~thq����	�|Xo������q�R��"�UlrY�n�M�kF:g�@!��L7�h��_s�����C����S�ʕ�������C��aƚ_M�����1���$n�y�KxR�:�E��SS;��=T79��{}�|Mҁ�,����:��yv�r?|3�������m[qwx+�a��rF��E�g;	L���5�$���v(f7�Ů�s�p�����']��#~r�t�v1���5 D���ާ�f����w��f��mҦ�׭��6�z&9�w��wS*g�q���b�,QQ;��92PGW�0`�8s�;�I1�jgʖ�6��ʂ�ټT�pbs�D�D��@������qf����,�Ʊ���?K��G�)�^Ғ-�\������M�X{%C�r��6'3�ǅ�d�juN������d���n
<^��ȧeǗ�� P�����q�c81�q<s�f���S���1'm�`�1�܊�"�	���TSń� ⾃�`מ����&z�v�����l��$���I�W��k�*����1��@yZΑH���Wia�g?7��{�x����J������[_��6MA"7��M}{�/���A�4�^��=kϰ��bz��z;gO��4��=���#0ëH�����k�]20���_a��D�g��u�
�7���ٙi���Ov�,5��<�@׸���S���U�2���D���ǔ�p��,S��^*f��n�C��Ȃ9w 3�q�M�/��Y�~��Cئ��J�9�4@��
���\���R��$͞��j�Tٯ��6Uv���h�P0�e�K��+��zUV��Kh��ǫ�I1tC�F+x��oҀr�l!�Gv;���2=�"��?GD��	8|���_<��%7x�|�.i��%.�PW���+��_��&�	��tlK�f��P�k���&��%uqɬ��Bwr��ࡕ���X�䅈�W� �N������o'��!W�Q:�=A,L��aG �*~#�,-���#M�Z;�D_��e�s�#
��|��k�Yl�B��|<�͍��?�[��om��JկWz���JT�����1�u��m���8���^+��3�|�^G�g����kM*�~�W�~��y۶Q
"C���[;^��6�3�H"St��E�d���
���ܹ�����8�/�R�n��������O�� r*�\��L��>�z���ZHjf�����ł�d:�/�?~�s���������#�Î޿~��^
���@�g*0��li�"�-�aA�:3�0�Z<v����g�qp�� f(%�#�7]�}��0}���A�k-L_D�Bآ���£Ѭ'�fn����]��:����h�UQ	��F����ż
�����v:xr�,�^_�r%Ī�2��PhÐ�a�QT�C�{ԧ��В�<��B}�r��a����vȌ�%�ͬ�iv�m�hE5#+E�(H{!��/��ص+�pߌ�k��s��d.�ʕ#]��S?"}\�1[�ֶ�=��ʢ/ʜ����&�QD'��&WnX}�x���>��0]�m�< �w��#��	F�;�藘�;�>��mZ�m?q�)������n���L�C�1B	��uN���{�B��� 1:��7���-����{�w`��e��~��X";�$Ə�����7��:�c�M���^dQk�a@V6p��r.�����"�&���_����%d0�:餪w#���\�O�jp��JټBc�y��l/{�(��wӆKpE�3���QbqV��u|)-���ܰ�� �*	n�*ͤ�;��o�� ����e)�JyF/M�U+�>�U�<��D�M[� ��.��4�՚$Ж�FK+@��]�S^�я
��*��ҵ��q���L����7ez�:�!��-(	����/�,���ը�蒍��{��I`7��h:@�r6τ��3P�q�n(t$p��<KL�`/� ��rä�~U/<�DW���Co:8|w���l�b9�D�±�xk�[�)��]�"�	��0�E�?�T����H���?�ڸ��(���Ip������������Fb���$f��B��,+@9�Xڕ���e��Ĵ{(��ϋ�ğ�+�i�s��F�U��g�>���+6l|Xe�TE�׊u&���>�n}H��G�mn����������lY7X�WNEͨ抌3W��^�.Zr�����a��Q��ވ���	�Py�����������"���5]�߉�n2^��hy�F��������i~��!�֦��lS�.}3<��p�;r��Q�-��'��qK�sV��:G-���er5^��s�g�C��j�0�Eg�q���hm���4�]���f���U"[܄w$�c XȄ=쀥Ό��6;b���F��;5nϻZSE/�I(C�쿋�}�Rr�$�~�5�>dv���K2�XN�![=�:кC&�^� ��>f�D�#B_�ǅ)9�&�k5�Y�������Z}W���&��rfW��'�����vP�Cs�󰙄7qL.ю���r���{+^̛9�;N\�1��>����nЋ��� �ے���u��6���#0��{G`����8��]��F��XX/��F�#Y�z���T�"�[�C���T���en祶�!�>�>w!}8�Oͬ�K8��G���5׿PG���0�;ˁ�^��Y��|D��tt� ��I?���7�D���K����_���3 ;#��B� ��ײy���������a�o+��k&e���U�'���Ŕ� � !�6��a��{�V��n�������o�Œ���C;|�$yr��}3��ے��Tp�!Y!�nD�㬼�;u�2��}��6�D�8pz#2`���iXl9?^��Ս�����c�1iGm�MK�Y��+�����P�p��
~r�9��sw�IqQ�`��c8�g��k騏�W��{�/l��w@�x�?� }�B�Qd���dg��w֭:�P�¾M����yX�¹�̗�>�-7��x��G���$�sa*��Dҿ�ߕ�7�ymq��>���O���~���!�Q&� �����׆��,�LoZ�h��}�����m#
N� �)v�����:hn�k��_�z�c��6,��^w~->T���k�3|,��=��k�2�w���u,v��^��a?J�N@���.
|y�H�(��x���1��d�v���	�D]5k�8�r���{-����~ �wJ�/ƍ��P��t>]0^�k�wS�[���4����E��Wj�#��qU���_�3H�)~td����4���<x�_��`ۻ����a���� N�/��a� ��o��>]z(��p3Km���c%�������Wd�ru��3���`��W�J`%�8Z��������d��4u��(�NV �2�q��|Wz�L�TkF ��ğ�.r�����|�y��=�-gǭ+��p�s�'��A#�(����w�y-�2�����̋�u�KGUF�_q�,�]ހ�?|�[��\΍��|����Լ2S���m^9W�0�f7��9+�g�$D��}z�(�E�6�2GB�c����D�KJb��d���{ ��n�}����׿ZL���%��c�3��� �X�*)U���At��u�h6Mh��4��Cs!������I7k��'%��Q��|��Z,�)�}��f+�{������q����nL��~�[���*��P�0ZY�������_����p%�V��x&W�X�P��Fhx�Q�j�6�9�ˀ�R^���>����|>�@�S,����C�'!# ���ފC�Z���y�G��^I��=��j�����#i6�3����g��������&y�����n�t�@e�k����>[6O���c"��Z���tFz�cR�7t��p$�k�	�LK��x�gAO5�����'!����mf��-��bf2�2�w��mȬ��gѻ�i��H�[�
��X��py�ز�rz�v���+5B������P�'q�~-�w���A�s�P*�La�?Ғ-U�-~:L!>���n���	"�D�f$o��2"'V҇@J�� �����)�s�t*��K����l�\GΞ~���˞��D��X��h��G�|�}gw�~��L,��KK��*�Rf��c��;Lbz� 	�"�[���W,����Ȭ��%�_2c���<��!��w}��_!�;s9��![o�4�yXg�O�[ٗ�G�5Χ��OU�zB�������9�+E��>��^e&��f ���+W�ϴ ��ȵ�^��V����J�(�=����'����i��r�q
�i�u���i���ᎊ�ٙQ͜�Ff`O����|s`� ����[����w� �+`کs�}6���!��e���w\�?�C�@j�:���D�ￅ���������ͳl9C�	���/ݐb�{п����w��x��o��:YD�"H&�E�HJ?SMq����D���#�4̿S��H!��
�(C���*H�
W#��?�##�1�TyS�v(�1S��%n�3��y��ߊ�#D0À��I �3��k�k���2�ϵ�����~����󌚨RwP*���}/�U��͈}��DEG�� ��:�*�APejR�?G��O�%ܝ�zU>"Qԅap,�`���s� J�)1i�a!�7��1�%P�=f����^!���x������$�܄״SlX*�qOP'ܛ�7�[A�[5� �Ў-sf�����f"��"hk��=?rb�@9��8���J��=���d��3W�ڙ=�L:{&\�shA��&�#���$���r��G���(���c�V��y�����)Y�P�Q�s�]3�N��'�9�_�6{�>kź�*����gㅗ��J��j���naN� KE�8!��KfkW���*y��:��l�)�����y���y!�'	f��6k�[�c\ys�Y�$��Ap�8|'EH���z� ����#O�&|����q#c̗�� l��<� ^���?���6D��f�$������6yG�Nzگ	�R����@�������i�hE�[*�B����y$Yh���.X�Yp��m{��MV�鷃膱}II�H�-�AH{�V��"S��yw)lo[!o���H��`��� �����u���0K03�
��'�+��%����q����Q��t?�������3�o`?���a��;�`!�>���a��=g=*������ߙ�c�۬��>�Z��}�͵���{�%Oh����lǷU5�����I���g�6��(��Ǐ�L�mjj~��$N����W2���~�#�i�f��+&��ⓐ_�u�Zu��tj�g�R�����]��\Lf���|�\u�;O���2m���/t㩤����-B8���l��r�O��=�� ;Yw��w߉��u|!��nmcZ���E��t�@ő�@cǊfs��?�I_Q&���_���BT�	\+><G8@���9�Q�]���<*w�D�v� ��^�T�#D5-�(�8�\4T�0����k�w
 ���ް��G��Λ��{�=ʬP��z3e�j/�\=���Ĕ��'�q"aҚ��}V@d�c�+��#K�A��\9ۦea] ��I_=4��
�����.$叶�mqN�/8�x&���`x��E6޼�&�ٚ>�0�!�=�/7�P�#P�hD�É��K{���ƅ�d7/�V��5�.ƗS�:�	+���|��Y�c�%Xyɇ��ĳ�d:J�P�0��������ߣ�81����c`Oj�*�W��:�#��>�q=|Jx�Zw^c����N�>
�C}�	�@��[�w�,o\���T�M�IP%zϝqm`��eC��O��MG�WTF�8�'���=m��;ֿ�x�z]����:D�I�/Q@��� �~�@"��TM�DP�4,}�\��zDTw�w�4gC?;�DK�}8P=>H��S7fL�����_L�H�㺗�a�N�q��8ky��s/���(�e/k!v���.��ueЯ��w]Mo5����S����_6<r�eM���~&U�
J@�I@��fw}ĸN���5L-Ť\��c;����5U(p֐4k�	�3�G���:������"PIz�]����\o������N�N�U��yw���q��^M�/�@a��k�e9��@��1Y�zz@�ҁ������	�+�UBj���#ƕ�1y#5"�ѭ$G�mX�Hо*�W)u��(�X�k'�s�2��_��� h�Ј�ʓġs_=���ύ��ЌQ=�|*������[�P���*�+?�q��1g�#������?S�?���7�
�}��^Xx�B����]$IS6�~�~��S�ݪޟ�?��C��N��N_c��f>@
Y���=����s����E9��o/@��wb�A�7��u"��}�j��?�ɹ�+�
HeR�P�~�(5�x��/��<���E����3S��F�&D��0&��G�d��F��S���W��o8�H�ڀ��[�t�;P~9sm�ȫ�F�_�6�jǝ��YW�nB��\F�[�����x�Ᏼ�%�< E�����#y����O�s �v׷��,���ɻRh+Nw��+������Hţc�}�+��i6,�.pE\��]�ݸ6_��q�Z"�W�Bj��W<W����l�����J;R'�,���b�*�����~zQ�Z<�z!��`����L��tI9�@\�h�:�0�4�ѤX����z��A��� �j��Io~#�*�����L�oY�a:��������.�K�� �DO�~����TCƂ����oU��<��-�:B
��v��iZ��Ιd�p����I*~�a0��Z����Փ��`�u6
��m-�������8 ���N@z���l��`��1�	
v�y�8�x����"-y�Tk�,���Bez��Y+%:��v��I�!������Tr���zFl8a5[��t��g{��"�ݹw���_Ú����%s�6C�R�(��lfDc�������>�l>���?�;L[��(x�7xC�w��]↕ܼ?P�E�\����U�02�j����1{��ry���ʝ���M5��涷o�`��A�:�i�l��y���`r�Җz`����62���|?�G���S���r�p����P��l��mb�j��0^�I ^R&���J,'Iy�z:9q�]]?��lph~��Äd��ML����U;�(��E����~���_��%���h:�5P8 �ˤ�@��X���BF�r�Y9}��ghc�o<��f��̠��6
� �}�$���e�Ђ��e�B��K�j��?� x�ƟnğC�>u(�e�b�U�a*����:��l�)Ԛ��Zި]�U�EЬW.��qz�B���!ί�̗:����jo�}��Ca�8���ֽ8u��0%�!�.���hB�n�o����ʱ�>����{�_�Έn7�G��w�r�i��G��$UN������}�#�e:���!�xs����\����e�2���J��"~):�Ď͉Q�����1K_7�lr�odkmy���z+FRa�餵��^?eҭ�!�s��w�֦��\���M��X�Õ�|g\��p���3xSmί]���HFa��l���W?!	ds�D��ꅑd�PeVS�V��3�x���@�Q���џ���[l@�e6%�-�Y�
ж����v�XEn�$S�P�'.�և�iHݦB�ޝw�^�� ���Y��18}�*��W�:2�!�S^m<ش�~SȮJ��5yGm]+�r���Vo�A/ ���"��"徭#��[��I�K���	 ژj��<����kޚ>���E^�?�7$��T��ժL�k�BHʎ�Y���]��-��&�N��E��Hʭ<:�юF.j˫�X���~��g,�*��9]�M��i>��Y#D�޲6�4��n�� �H���� �95��딒��+X"p8/��Ҫ?�QP��e����������ҍ4-����M���)�E�ځ���g���I�PS�L���2I�2�D���'΀�� d���OZˍy)��\���f������ut����TQ�� �-.�ǐ�X_Q�ߴ)��c<���P��jVƸ%?����K3�����B�aqH��'�㔓U ���r�H$�5�^��A[ =3K<�v}:d��_��茙�FlƋ�5;-�>�;�K��J�hIc��Jk��Z��6���*`2��_#��<!/��#�.�����)d[��[�J���pJ�ym�~|�A�tK��);����ýg�qEKG\Jl���p�If��ꤕm\mF�|����Dꢴ����ͼR�{����bb�k��:��_�{���P�̇�� [WZ+'Ơ��?F��h��,�T�˨
������:_�s(��V[F��ȇZ�@��4���!eѪ�,���/�H�X�@}����.��r��V�ہn�GRl� �j�����襦��*���x�ﷃb_:f�'��1�5y����>�6 ?��b8OQr�$��h�ᾪ�ϙ(t�����W+w�,/d�e����%��Z���dZhm8
]��?o�����.0���\9o�c���͔R�����p��7��s�zoq�-�	�Q��.m���̳h����qHsnY�Hv}*�g_��DA����n��C�7_�ZJ�j�7o����X�!�@/\�ry��с��w���<����L�0X��������J\��$:R�и�F�:Qqvb���#�`�l���_�8�X��y�0YD#UiO9w����Z��ݜ�|��Ȁtz��Q�-�x3�n �GwqW(h��]�T�0e��i)r���c����ed��	���gS��l�y���5E�3FV��E�b�[�N]ɇdf���̙š��G��(���`!�GDF��q�z�)B_�)w�̲����;��j4�!ߣ�g`m�G޼�,�n{,d�VjͣM�X�1�44WmP�e�
V�G�xD;Q���ZW˨�۬�w2x{[���ٗ\Ϝ��_�՞ύ0-�5X��Z�ԭh��̘�ןU �'s)�6'�4|�Hw��r�r��t�ǟ~T8��?���w�qX�����&�eR�Ȱ+��I�akZ�
��nэ7�W&�CbG�IƄM���\����+��-%o�k=�΅�|�	����L��mo2�"�(ZM�/�Ӌ!�O�8t���$Y|�/;���:r2����H��1�\C���u�E��L!���/Po�|~���m��B�i_*d�f��-�N�c �J���|u˔��ۦ���V�<�@G��5��&r����<��mq�#��^x_��)I�2����z9	��7�7P,�z�u�yx�t�Q�6�gr�qB=L���% U�,�,���:�:�O���՜_���O$��bK=���M$I�k9i�;0b"���7������?���+�Z��J�6����r�5��w+l<�>_�T��lJn�qn�-}�\��E�G���ƍ��J%�c���H�0RJ��5_�c �WY#<�؀�pg���|Ii���61͸&#��tC����߳�u���g��?�*��mw7���II�/���\���j֯
³����Y�oBP�;��ބ��E2 ,E@�2./��|/t���N��<`�*	b��Ś2z�l��8�$u(�P71u�/Qj�?z�=��Ӭ�����tk �UX�oӁ�����,Ib���P=DF�"Xt��FTuE��`�rt{�K6_�[{��}��iZ	 1�v�|����+=l~�jv����ߔ_	�m��2g���eI����Y
%ӥar�yK��	0���zzh��(2�l��*�	���ĥ���+uأhz���+8���
I�#!�`�$#�_��@�{��y�f�j#P"z�%��OF�SO2M?�y�J������5��N�N�(�ϳ� $�U�X�d�\W��b��P��I}����֔���wl�	�!�f������f:���t����D(Fܰ wW��窬�gs5�,	�^�Z����f���;к�o�[�擇a,��Q=�2�Wc��<��M����;%�	�Y�,���	ލ�O�.���;�΍Kv&J���m<�wN�1E)��̏���J����t)��(e�{tqZ�N*XI�B;�:J��z��± �D����1��K�;p�ƆK��y?���"��'�(�-w�~���lX~�|���Ȓ�e��������(r9 4�d)�Mp���;L���az�&~]�Ҟz�!�������Ggj=���7n�|a&�~بǉ�<38��$�Aǭo\.%��u^iW��JP#?}9`��ԝ�dF�[��6��@�Z3�{\Py9�@�7jX-꫋R��ͅ)��H84�T��������c�-L� ,#?F7��)���T�X�J���"��l�~uj��{�a��D�Ď��fŔ��n@��9Xc��.Ǟ��,��~U>���)�Tр�aSʜkډ���[��=��i� ��.ǧ��A��|W��TI&��-+��+ ��Y�%��U�TT�LЁ�+���x���(������B�2@2��-ǈ��[Bp�N�q͑�������M�Ӂ��/�@��qD�_%�K��T"}
��G���I��ef�j�Xyw}i��nW��A�,mS�o��l��L�o4�qy�Dp	�[��ҭ|���ˁ�'�ߦ�K.�M�?�����WC��!p8�D�9�[�p��!j������]i�7���C�����Y�D<�7���Z� ! �J��ʂ銒��^:��x�&eǚN]��:+/g�{bȶ� �mL#m��}z�o_!����D�/t��*�����s+ˤV���'/&�V�_K�55�ej��H|/[d�Yz{��ǝ�[qv,*#���h6K˗��B3�؆�^���R߿T�[��홳���.���������A>ws$��eW@r������#YPs�u���Un"���y��~��.�>6x�66��4��<�S^��R�!�����f�����F�&��J�k�o�|����9���G�g�c���yΑ	Hf���QH�������K�/���q���M�w��� ����r���Se��@DX�x��aH)�դ��JST+}`ɸ�W�oʪ9�L�:�Mq9a��猴��4@|�Z��[�W���A,��j�.J�����x6��{�X��y�x+�A��-�צ�iVB�ؑ��QC5k[��z��"@�����n׌_P�����stPu�˔�����o(u P%Ĕn�0��nC��D�#����Q>�'�V?�%o���/a�:�JX535��j�ؽ ��y
�=�����j��h�R���t�o���J�P]��}���<)	�[Y@NU�� ߕ5Kz�|�2��O�'O&]};�}�ˏ�����}īE6�,���O�Y *X�o�vx�2��h�O��V|2���%Bշ����``����N9�`#Q ��u�j�Ġ��tDK&M8���T:=)�	J�|X�VcF�^YGʂ_({� d4	�3(e�����$Gʩ��QI��1)yUG�GT�x�� u��9U��e*K���6P�w����C>��Pש��ֹ�4mg�'V��.y�4�L#�� R*<c���g�y��d=G�������m�fږ��Ҭ�B:8E�+�5�ì�G������aQmo���
�������H�P*�%1t(�!C����HÀC��]����0=��3�ts�&�����y�X{��{����؁Q idpw�	z*�O-f�S믷x�N̧��$���G�3��2|6j�z���_	ٛ��O^5�4��R�R��L�s�2�B�������V��d�y/eB���Ǚ��0�j$ ��ar��](�]�}�~]A]6|xz�I��m��?���~گ�ˣ����lbS��i�ʗ0�A�!Rm����<A4��4Pwf�
D�}�_�K^�0h/-�v&���d���[�̉�6�"��B�']��2�����[4U�%�H�u]�GRԵq��A[�H�φ��a�a�^mF��ۏ&����؁iƖ����wo���#7Mҥ�ŕ�;^r�M��0�[�^��ٟf�/�!�(ls�[���o�V�����Y��H�o��.zo}�2	�d��<���ʙrI�^�V��^ۢ�ٌWA�e�i#o�԰Z�ln".�	6Ԓ���hu���˚�$�ԯ������pA�ű�v�t�v~���m`�!,ۊz� N�f������6t~;FK�yH���÷�M�|�Ӌ�b��Y�Ǽ�_�_�)�D�Q`*�^�9�~n��:"ۡ9���z Ù -��I���s�y/n���1�*wt�,��V�q7��(7��S@�GF<~ ���8NV��@Y
�k6�������1�2+��"���MnWj��d�y\��tu}�5�N+�}C4�7.|~�G��i�2��^���)�e��2�%��!�֦�S /B[Hxmw�4z(�K+�!VI��X�;O]�~��4��N����������9Z�ؒ��hni
a����y�r]������B+����49�Ia���`����n&�-��ߞ�ˏQ��H1�tv�A9��/̄*4�ī�R��wT��ր�\ �e1䇾~����͏�5�3&:2�+C��LVYLĞBY�v��=d��Z�_S�z�\��Q^a�� *}��Gy�S5�ꦵ�e��jZ
C]�{��N����M�7jq:,���
v�g[Xn�s��)�h �I��j�.PIb�-G��L����>�Df7�q'�v��.KV������K�#�Z ��,��k7�>�g{K�����$@�P3��e�vuq���<��HF&�^.x��&@K�� �| G�A�-�`��'t�r���)��3�c��9=����:M&<a����ne����'a^KZ�4wFs��p���8���%TA@^�Ҁ&��-8�fG\�I ��
]W�p�V����}<�8a�U�-�w�6Lkƛ�	� ��B���&�]
~�i5'y�!ħ�B�4f� s}�� }�&��ƀ]�|��Z~���7�qZ�o.xF�1woߒ�A��'GH#����
v�r��:��,�A�'�e�?CE֒�����׮���xK�bru�h��T1��a���U����w\�!Y/%lB��\fn�ӂY���N8�QhҲ���9J�n%-��?��k2�W5� ʢ|�#��\Ѽ$�B���̈%��C�xԜV�+]��`x@P��ߊ&���)����C6a��
I^�
����	}�#�B�&��s7�Pn������a�ҩ�O��jn���N���{�B���m`��}�����S{���2��l�!ť�U�U gw��t$���&&A�?"��,���P�2�KAN~d��������֖�T�S�-��)�����#�ՁB<�����ԉ�B��N�a�k�Q�l�2���n��cy����\M�K�(����їB�b����S��Yx���o��IY���y�\��|m�Cl�;�Jæ�&���:��Ws�/�ȝǣ��tBū��1}�o�����@L(0G:Nn���3A�e�)�,1�n�.G2��  ���c.�"��b]��Zo�[��K�¥p���V/��J)e�(�~T���j������rW�,�u.�v���fY�qS��^Ļ�J��V����w�L�w���:g]!�!�d�zcg-�	��ڸRs4!X���ZX�FRy�UT�����s�̭�N ���tY� �:�3�8��F2��������m�x�=�5e�K�gk.�@Bgj=5���c�Ϧ�����d~�Q�\Ϭx��}%1yݔ#��>�e��jp�i�a���^�~�i�{�@��n�]�UPѯ���X���6'�f:\����NL��M�|&�Jt]˾��2</$��s��AH���ڳ������r�O)���@ql���?j �7�i+ii�6b�݈��ޤ���i�f}f���~�UſU>�ŷ�9�yF���] ����h�0�	�NE�s�ګ�L֤��A.M���i�"�x�>u�0����*=�T��N���4������a?(�
� �ycQ���|�^�q#�d�GZ_2#���DA�ƫi,j��	��#��8?l������X��BVY��/�~͉ʿm�������ͺ��m韋���}��<�z���!���Z߹)���^���(���B{����c|��D���_���$�u�`�hG��eD���XwZ�|��4��I�e9����$�M�����F�W���67O ��=�O�=6��Lqu�8��㬈"!�h.��nd��O dO�U-�4�z�}ˑڟX�)�k�D��]��*>Y�َ�J�����G6���aUd#w%����3��+G����e]����u�׳
�{�� 7)j�D.�D+\zטl7ݱ�a#e��=Z(gV��Ί���j!�]	�NG���8)����U9�t/'`O!���D��B�L�J����R�Cf-~�qC��^��5ʌp` ���C�]M�����3�}��5����'C�F+��n�����8���V��p�B�\{�rX[3.�b�$�{L@�!Kyf8C����b#����G��zHW�)��!�m7������Л��-^ޡV^�܁��ߙ��o�s�N��$��ywL�D  ���!HTTs'�����m�f���̂A˫b8�� �g~�\�j��	�Η��̔9t"^�lb�MJ��1��v�P�+���>��bo�:��~&���븍@4R� %�Fe�̌/.agC��^d�g둺*���M.��䣕�4T����6�:e�<O�>r�{�ސh��<���K��ۣ��P���2�-SJ����Z���ʵ��Ri�$��^��^���K��C���"G�,�O`�ˀ��6�g����ܫQ2�c�o�|�s�X�b\<�m���Ya�~]Tg�coo�%z��	��LW"��QP�ȿ=�f��;(ߠ�JF�v�?��
2�/<��_ͬ�F #V�?���s�����C���n8f]��
}����\,R�O���eɯ/e��G�~�2�s����o��'pO��F�����]��"%'�\��P`�K�'����O�����Lhh�� ��R�u�JcB��r��8 ![�g��{�<F+@��r��S�-}ju�~��ZWL���v�fv�Vv��܋�ɻ`C෠�<Ʒ��d7����>��d�;-��NH���ޅ&}�;z ������2�����Q��30K�JEPb��Ml�����~e��٠��/��m�T9��$_��366gJ+��M�7��!��(�꽅&9����O�,�MK��A���_�zˢC�@m��Z�fue�Is��}qң߃Ҭ�H�2�c�5/:{��t��˗38�0V�~|�Y>t/�ƣR��mr�8szm���C�0���w`\]��:t�K���7d� pf�ds��tĝ&������d�7( kݰ��i�J:�}�.�W�+���p B �<�(��}u}j�O���^�U�Y���=�l�����|W,t�K�#�`� C1�E_��B[u�6s.��uN���'/��S�h�0�{#%i��2;
Y%\Ԝ�O��p�x�&���J�ji��	�_��X���X�dU̯{�;Py����	+����,2��VP�Q/@�P4��K�i�C�̡���{���� ���I*�뜆0i��-DQ+��b�4$0���2����t���^��ɔ�Gv(�c��+�3õ �9c��̥1]�+��~f,�4w^�|+%�ꐩV��V"�0��]T�Q�R��o(�<i��6z���� Z�	��B��?������^����1�GOw��϶b���o�ӿ��1�����W��v�o��dO���R��V��]��Lv�$�����˶C�+K/���[W�ZP���c�Ĺr�)�%��\}~�	K�L�޷�/��� Ny֩O��Fٕ3-�T�vSV�i����Y�f��_w�)��*e�����
o�THpg�D?��b
o6dog�\\�e�G��~5�^^�H���P3����,C~��#+��2���������:ɺ���#���"�TF[��)��HP�MP�Q��G�c�P5�]XGe�xFtZ4����R�K�URs�M<���#�_AK�4�Y���Ĭ�,��5���g�}65)�����
�[ϗ���������ul�;
.ɯS m�P��vW��OqL�z��e����!��≯�s~�P���R?<U �/�e��Zݲ+2@�\b��=�����}��xֿ�g�C�/�%Z86?h�9i{2S��BjB��D�=�����J�̱y�J��Nz[p#4��-L�&�����v��sr����6��,�owj�F��c�X��D�?�Y'��.�{�����uc����r���h�΍�U�)D����=�@�.�z���*�#+zMK4�T�b��9����Q�V��By��Mu1��k+dLŴ��X���_E�Od��ǕCy�|�`hbTȧw����N�����@;㻔�3�;�P�e��
��WE� ��w��٦&�V ��鉫9�b�i�h�����--�qG���M�T��r��bZO�Q���fY����n�) ~S����������c��_#�̑��ue@�X1�`8!��mfjЙ����8bAjUW�@L��n����чh�H	��aъ �m��Η��ű[t� ��5]����	�p�oi��0�(>�Y�M>�Ө&�>~�Tǆ���U�~XR��0�A!׏`"�Y����u�Ǧ(��Զ�,���6_�(�ң�>�_ #��L[M�{�U֣�Os��]qͷ�̜�^ϐE9-��.D�+8�b��`[�r�� 5�xB���|�3�|�9��]�}�V��x�-����ŉ�&ɂ��r,��-zѾ�./��di"�L�#�`cg&c�^���w8�=�?�I}6U�&*E��M���C�<Ccm3'��Y����3�a�#��O�󴓀�&�Ԕ@! �dX�|'8mf�[����C�$�Z~��^lu��S�p���O�����n,B�	�)RF l��F��V�4�B�@��wSi�^WL۪��g��&F�_��<>�[i�4Ԙ�R|ͣ��i,��G�]�V�� ��8�#��2���]j(��4장@3Ⱦ��I`w��ˊ�*��z����I�n�^���HF4�W�xU�m���G�N�mH�V��#ˮ�m�7\�N�Z��UZ�堲SQ���o��D6��c%�nS F�!vǹ��W��k��39i	o�O�6����R��H2^�{�1t)$�������{�!^�9��F��~u�*hw���ж7n���"�!��iX���`��f���`���uh��@�����u�j��-՘I��݋�����h��j���puR(�cT���!�|�r�:Q�E����}UX���`�y�{w8�f߈�!���X��2�.K��x×>� �q`ˑ�莱�>��7�N����܈�	���~p������i`�����Z��J��w"I�W�ࡀ�u�EqY��=)����'%%�[��syj���|����X�N���
׫�I����gfN�%Aܐ��� �0Nu�~������U����f[� �}D�eok��2��K�5��g��:lB\?�x�W]f랩{���H]ڪ�k�c^�0~�%Cۥtj�+S� Ͽ# �>0O�%�W�5��6�K<�!p��=�e�M��ʹ6����jn�{���RG%~�ٯv�D��\�x��?܄^��Ǧ���#T@8�!���=�+��VK4��WZ�yRe �R#�����������V�!.�ǽ�	��0D��ec�pC�@K��bƋ|I�	�D�*����[h ��r�z�*!�;Җ:Z#Ӽ�?�F���c��5?�U�{\q����!���;��@~�b9@���*���{qz���$>7�Yxt��'%�9:�&LP�x{�w�Iі�n��ۆ'�VН9%tߤj�=�yϭ�h��������P_=~c8�D>JV|yW�։�����z�`��p�;�k��\�%��>ư����rVݞN�+
�T�ļ�tR�x��և�Ȩ �����%�2��Wc���c�CR 7�hH�|��͢sb���!�>H�s��/Y�'5k�F>��<�{���ދ'���N�^ށ�J�?��9(ޏw¥��0Fڋ� �a-f�?�q�F��t|楓95���{U��>�T/V���c�7��ũݍjY�����3�W�2�� �Ats�&Y�$������ڔ�Iv�NO���L\Sɵ���5⧃O��񉱭�n���]���y�v)T���	�&��y���	8�/u]&>a������3tC�Pc��л��M3v�1��������Q�^���)�K����cܞo���z�f�{�񿮷��N��^�[�~ ��j������ﺇ<ZR��ƨQJ����!��/�W���$�X|uWu܉���h7��+��o# ��6��C�90n��۴>����̲<�צ�����lqf8 
���(3����M�2��w�O:��nf�[�WȢP:9�lT��d~�Z��];�4��H���g .ue|g�r��NC�d�"��r74#7��b��U[�\ݺ�Hw�Q��a�l �@��ۂSȬ='���y�����f~eO�o�x����R����ѧAV���,�ŽuJ��t���e�)��U])f������u�͈W����x�~&��-|�
_�b�L�Ņ�ҡl��Θ��Ǳ���^���6s±����2�����/;�C�2ϛ�w�.tM&�M)UJ��m�ـ�v��F �}n��*(��F��9/��l5&99�3z��gf�nf��
2zkV̜��zIJB�BT�!�N8���*��.�n��'WZ3C ���봛��N(G��m��3K�X�#�P��_�<v&~S��G�hD��|�i�F[X]	-yqz�\jȣ7�p�b�zg��(�gA�K�u%�F�:g�QjϞ�<�����{�kh�VZ:���{\~��e�27݋�;�|�#;��Y!YA?�M��=Ų��I��!���������f_��!0�7�Wk��|z��lPh�_����+T�i��
�����ƢZ̩5.ɿ���z�r��G㖠�Q��W`�`��9O��w�_���]�R�UwKF��ɢ��	C��b�����ː�X%�W�bʉ,
_����o͈�
rg6�}8��������}͊��e�fH�H3
:7|3>V�4>���YW��i�5?;2��J*�&~BC�5�н����%�k1J~�9:Y$�8��Rʾ�j�B�'7�f�?F�狚w��)�|1�x[����^�y�hN����}h��U�D��1�,�j�T����{�v@�0y���R�7��P�w7~���o����f��  Qu�ˋ�����2��G���I�	A�wt�#�U�B�6��\��w	�^d>�M����n�����я[?�3�˖�Q��ne�Ǜծ��P�R��K��F��[�M!�{�sY�B/K�G\s�եj�LʄYѳcY$����yC�G�������(�>q���(�ݩ�6��� d�~˞'��T3g�m�N�dP�����z[�G�Yxk*�x�̚�ɡ����S���G��V�l)�o����aދ�	Ix̀�=g\
@$Nh���t:�� ��q���l�����I'��.>�3RIc�t�c_���5�u�����Sf�ben��Bǔ?�"����ٖ�[�mv�x]}�T���P�~�i� �G�u���]</�υӦ�����
���^q>��ƪ�}���Q�)е���L��-�����)��%�M�͈��Y@(���B��3��d����)F�H� �g${���'s���`"z�����v���߾��M�{VKud�>͈ ���y�.Kq�COE1t�'.���Y�:���ʪ��2u��ZJ�랛 l��HhU�_yZ}{aV)�QS��%L:l��}� <G�*�P�Ua���S�'��(o�uu��f�i�V�� �mo5�b��f/��Z�ރ�p��Vwk�1�?����az��08�E����g
v�*�ܤt�L�V2�¨�pǴ�d?-����-�F<� o�j ���V�6g��mP�x7�J����V�Ek��d��hN��*�8��
��^8~���@H�s��ש�b��9>z@�CL5�^����W�~!���^��7`Πl)s�#�Dl�7��P�&TC�5������Ik���\�4��|Z��{%�zϹI�4U�/W������}(��p�__����rfW^}��k����m��*M�ӻ�����ף���a��E豞��D����q#8�h��Z�ء�Be"h���N4|H2���<��n�Ѣ�uW���0���GS�
��yA�`Cs3�!��X�h@Y����ў84�=����P
9���ʃ!�%�ҺF1��$z<����LT���b1�Ai�ww��)L^;���-�}RQ��6��gU�c�i�;����'A��v|�����a���^=Cg��i_C(�@�%xp�7�S�D����З�W<�N�R+)֬J�q2t�S|-9 �m�r54��RS���a�m�	�*�/ � ��:9s���&?m`��W��5z)�{�`���۾�U��;*�L�~��u�?�U�D�{���F�;���
��@�b���Ǒ�)�)�.��?�ԓc����U�c Y�@Y�!~�4Im� ĵJRD�u�;g� Z����e�~W�1�b��e4�y��P��F!_�g��]y��B��	�}�A��:��UV={s:�&�i5;����Ƿ�՚��3��KGpl�kT.fD�^I��s�4O�~�TMjݲ�T֩�fU{{�Cy��s���#��H��m���e�#a���Y�B�)gK,�
}�3�-i:s��?�Z�)���$]���T����0�It-�`gKY�G�y�'���o�8�WU����u��	���,{����}�R�
��+8����祖`��fbD�&Qj^'�0��O�$��V�wr�t�γ�>��<|���ҵ����&S� ��bBcT������P��c��Ϩƛ����yف쁰��g��S�����~�N3+�"c�U`e��X�T��ZP����!i+���F��3�����i<~�ú�f���
��f�������w�=�g̇/����9�����.�)��
F/j&CS	 ̀���*3e�����әF	F����'�4C}��e�-+q[�%ko���~T Q�d#����|�@g*� -m0����&�&L���'\hGƍ+>�6D�_��Rי���W��rnm�O�i��v�q`��}�.�f���#��/m�x��p$ɫOǛn6�ě��o��sRvk+�=���gUQA4�^����9��ʶ�^i�^�ɗ-�\�h$(������-�`��"����~���L�.�!f~�Z�"v}}X?(�<�Q_O��)�\���ݲy&,�Cb��gߵ���vwݗ��S�����wl�;q?P�;+��((ʘW�B��x8�Qg��*���y�s�� ��3#���#���g��T+��9��Ļ� a+�w�!_�B�đ������]2�W�[�)ٱ��3~�w�V���s.np[dX��9���s��k�ЛdT�/�i�t�垱�2�����b[�)�I���y�aO�]��'o�w���ν�3�U�P'
k���1>�T��I��$�kt7�5qD�9T_��"{���S��)�OΝ�;�(����Q�$����zr�i?sG�!����k�1&�#Bb��t2���n�NF�笖qs]~3d0���Ob�XFB��s)�?��0]�V�w���2��b�Xv\�z��fl_�vyxB�����uF�d-���e�߃��~F�R>ۑ8��-}>^��x�� a�3�K!>�n���l��>�?�������uwy-䑢�T7���5�-�����x㧲�Ũ�a>���l��QC��R]Ԏks��bSS|�%�;� ~�`5Q��ڀ8MF���+ȟ(���k�J�q�_���P7�ӫ8�@�*R}���Q��aɝ��!��]�,i6O>�*Vp�V��3�x�i����^Μ围�.�P��	Q^�o!V�=����yJ[�pL��_�<���\�:�Uq��0��t[7@6�!��ӧ^a���8���\��d�i���J��E3��x3��R@��fwѴ%x���e�MĢ�ZDD��IxaB�G_Yڤ� :}�e�:����k{�x��g%x����>
Y�����+Q�;��|�����';���)��=r�'����`����y
��E�/�Ҹ˩J�2%�vIUe�l��ݙ�ՙu�7,F��p���,z.�	@&�
]>�C���Y�>_��_�����j�9�TDB2�7X��܊�[<�Ә~�����6~�A�bﺇ�jW>�B��wY��f��ήoU�E>��~$O�.����������Vm� �ꥼT�Y������`�O�3=��?u�9Ҍ�q��3�#�W����B�q,'x��#�Z�	��r+0���ɣY��nzR&X�"/޻�J�?s���%'To��yI��GOG�4�e��5�>U�I�8-/��L�d[4G���|��S�8A�Cl4��2��?8[��z�.�dk<��\q�{+D|�Q��F3�v��ؾy|9�z�\"d�n=穦��}y���/=�w�VM~�bQ`=^ �g� x�[!&9���]d����x�1�k;���Ǚ�fԥ�h{o|�����Y�Jc�/�9[Ѳn��O�k?��x��������V�&ݖp���-�+��3���8q�{*�3;�$�M�,��-��BH�P	/�Ԩ�����+�@����Z���H�s�y�b���t����kް��#��=�.�)�.��s���Jq"�o���z}*J�����ɴ�r�����g��DL�կ���<
v1��G���(4�J�7~�6�Uᱫm�DV�=�AoN���Y�	��ҳ��s��ci��+g�6�����Ta�t�xU��e���T��S@�֓�a��8AhN{����d|�sᆎ�.C{U5����E�
�w��,	���wl(ޭ�N�۾#����	NhҡT�c�����S���/īd���'K�<ݕbA#0̶�Iȁ�<w��A���6����. �'x����}*��?ӕ8�����b.���
�Vwv�2sH|vɼد�y{�pp��c_�_�L��i���qY������-������lޤ�L���7�0鉳	� ~�дl�f�y���v��A���-k�B3h�7T'�}�+���9�^���gH,7n0+��O.�����u��(5/�� ~�g�#���3onz�p�}����;U�^/��:mHO9��� c߰J�A�"1:p�Mɷ��c����7�����k�������q-
_!��L�&&�,e,����� <8��KjCݕ���t����h\���4/��k�R۪��v��(�����ȗ�ڴ;0��V��b��!�\b�^�}y�m�W�oQ�B~����C����r����st��*7����6, \R���)��c6#�ރhʢCC�����GǴ�csE�=f�g�k��x���z��+ռٝ\:�������3$���a���P�k�)txZw�g]?2	��3m���>(�=�K��VtZ?Na��Ȳ�(�\�,��{V��) ��?g�9˦L�b��w[T~���*KI��;����/&�� ��5���=֯0yI�G�rENG@e0���Z,�`������	�ힵ�*��Z� ���8{���I���ٸ�myNm�HCo�^&��ħ�S>|��V�X�]�WQ��*��Sz�/je���U3XG]���6��3ξ�zh����X�):���egN�݂�`�*P6K'뼼]�ojj�G���5�*ϰ�G����i-��ʧ�w��ۂP�}���K�To�0Y�*���<��1s����(�'�Ε���j�r����x�y{��|�P�{�)���W��?��U���c������ک��'s��O�_�p���-挙Q�����8�Ib��J��)�e�߭���!�WS��$����*����0m2�N��o�`7l�`����⸘�������Ni�������+1J��vk*��̼�͏V�K��m�������b����L��u�Y�* ���h�X;_9�l&,��U���%��Ηm`,����ո�y�!�9�p�O�̬��J.`����sX	f��7P�F%e���՞��?n�*���ˍH��/e��a{�W70�4���y"j��c�j�*�������&S��*��l�NOg���~�����@L�Z���>cMU~�{�~a�2d~8�
Ux�n>O>I�<����<�:V=;�s��N� �M��6��ױ.�uF<H��n��ǯ�;?|���T�P!�[��g�nh������n�����[�sc"������;*W���w��/њ�ꦒ$XSb0��7W�,A�Rh�jr�>�f(PssH�#<�n�s�M�ۆ%F���P�p�^[*p.��Y�f�|�Yǲ7���w#�H�e�CaŪg(�A��X޼���r���n,�n����7փ?3 �R{�t]�.*�kY�Q^��o~+�5���O=��2o����x+;���}�j����bb�s��\�lw"g��{�y�h�=o`��I˫ę+��N�rܽ�$qp�D���+`o�Ϥ,T��_K,�Q[��&�Zhk��L����,$YC����q�}>�j
i4���ܝ����duT�he�T��rM_5���XG��U�k�-2��W� ���)�fę�j������� ��
Y��<�������@��4����9�֗��W�_��K�>u8�'�3������K ���ف����9�r@��9X&ӴT�Z¹F1-�r��*#{�t���~��>�7�^�]X��}�^�ft��v�
�� Qܹ)��5���p&T���uY�9oE��a�Z@VB��"U.�)Ǒv���ږ2��!+-�^DS"dvIӌ�O�� �ӛ��xš\�z���Tl+[���\)��S�|<X��&M���1P��C�W�oH|�Kq�?�˨S�T�gWL�Iv���K��~���!��#`�#9��ڣ��U���W�ߞ@}�
 �'�95�/RT1-�T?ɠ�PLo��r�$�ݮ����x��K��o��A�
r���/v�&[�]{��ej��"3��8����x�Zo�ᔹ�ݝ����wǷ*u�7�I��F%��@�2z��dؑ4c��͊C\ ���E��6FG�M�y��R/u�o6��pה	�w�,�����<�@R91\5����ũa�җ�T�}pwTrBP��1�0	K�N���=y�!>����X_�a���������_���D�7�ݮp�P[�*C�@I�?/�Hx̲\[�E�$N���#O��_|���}���=�R��y�xU�Pj��Kl��ȷ�nc|�]kpl�:u�y$xu�X�mw!�S@�qj�n�,�ې бa�z��׮�%��3�����a�/׍>D�������+�o�<;z��ߜ���Q�L�/Qj�8'���D�K�kpT�� .�Q;���䘦��ò������)��C	_�(��ٸT��:��`���D҂E��_���гT�2�MI���B�m{T
M_|׺�������\|X�K�J�����Kfu�ҍ�3X��]�ft�@�����w�ߟ2��u~��*�
,.p�qM��愾&!`�F�� ܢ���t@>�s��/D�{�Fv�E�v��n�8!�tͪX�!!��&M^����L�8W<�pI�#��bi6��
Qh�B-�X�k2T��3�'�Q����$8F]y(�ۀ�1H1ͭ3���o�!�:�%X���Μ�+F�O.��*g����Oe����0�T��0�xM- A�5hk$��� ~�Q/>��e�2*�k ��[��(�����03TW��m��4�C���Q
]PNN}gO�$��q%�(�!B�X�$\n�y^���`�m!��	�Cy��?5N@Xn��$�� p�
�k��7O�I7�*fz|f`�?!h�}�p��N���J�(e�qTڳ�J���Y��DH��@�(K�����^1>20d����R��*�̱j' �rJw�c�X���!��\�<���Y��h^΄tm�0�[5�
�楗��ۃ�EoD�����֮�hcL\bv��殤���2�Ju���Y=��y ;�p��Nr�jMu��>u�g�Ie~��4�T��#�S�L�3G��os��)���:�}ew``f�u3@���kbU���-�(�m����v:�s�;'�
�K�p��v-��.^�G�݊����Fc��S��������(���yL'��oGX[Z�W�|t�B���ռ$2��5<�GW�S';����϶ū���'f�Z���J�ιI9_�,���fP��GH�s��9U��t����e� Zd�$VT,]����j�t��*�J�5�w�QE rԑ�k]��BX�K�vf����[%�W�9[?%|�>�B��!��q"���.g0B�qJ&98�s2]L=�O��(�i���=q�~W0��������6�����'vǻ����cz% �RZ�k�;��M�FU�P:�8V_�nj,o��w!&(����6�l�����IFˍ�8g�&S�u����ƴ$au]�E`���%��o�p�GU���H�m5�lz<�B���@�uJW5�i�┎_�Tbl�����]@r���Ϭ�����F?���׆Yo����N59Y��\��w�[��(�2O�Tx�_ơ̈̄��$&�ь&���ONZ�O�/mpC�:)�Y�Y�=&�ה�OҌ��:��ڍ]|h�1��)=E��ӳ�俇uf@��*�H�
0���(���D�A���I��cɬ�P�䊮W �	q�,OxVH����;��o�o�7it�y;ߙ1���mZܷ�D;�0��"%ǫ�U�&,�W� Bм��6*�3k�6������2�	�ɒ����٪�C��+���$�(�<:�oAm��I��8~#vG?=Fu<tzK�yP؟����Z�&҆F�RsX�ICf:��MOj�����Go�.�y�Mq�4D�x ���d�$<�vrGT6��X�:01UbY�=L��Dx�tCf�1��xĲ.ˌ�Vl=�`Um����?rw��(��vE��d�Lk�J1�A��pcbi�;�lّ����W�؁7��7��e�������7�~�k�_�t�����Oy��%��"���}Ph�k��T������F>;��M����נ^0"ȟ2�`ŗN�syW�&ho%hL�L�-�U��HUa>>n�D�LT6x�E�k�ߔ��3~�U~1C�`�� `�����;��j~yHl;L)�5R��o��"���˵��!!-G��{,,��y��颫�0N�j��sܾ�s���5�V������"�~����ԙ�,�Q(��J�$��G�ޕ5�h�驜�)r�1r�ؔ�pu�-���l�)G���䭺[Mv�1J[j�`t~r��#3�C:��w�g�>�۟��Lb�O�=��R#���`.��Ӯ�tN�EB�
'KV1F��5~��I$��z'�^��Y��	�x�"��y��"o%��Nn���#"����A�?fQ��c��eg�>���iV���?����.?�2�����TFV�-�T4�J-��	<���^i#	}�Q���_ڑCN������Xtj&�l\ƫsR�8Hn���_�l�罐�O�ήdψ�_��S5_���[�h��Z�ƹ��D�ц���zi����$��0q��'�W���P\�(�JE��N�������>���D��Bi!F^�>�h�/F�V&e�63C{f���ҁc��C�Y����?z���<LE�V}�����ap`���VŋtT����"]�#�U,��SGM�$r#J��KwM���4Ę���%Z�a^V1,���������K���bM�lq�OX�v�����_�↷�2��	����ρ1aؘ������'��9j�o_q�o�h�>ۑ��_�G�t����w$��ͧj��9����yf���6k-�h2��L�`��E�·nppK�kze�VyN�0�����	DrּE'�,Y��s����=V�n#wd�tH��ו��(���Ω}��S~����_���̴�@�"�[��+�}�R�D )��y@�u��؅\�*�WP��Z����߯l���wJ�lG��&4$[�!X��XR�"E�������L��H-��u����,��-���߃@�0&�9T؎8��������A���!Ln�Bd�0}�S/�4�8�N�&�AaX�P7Ű��U=�"�o���5��Y?��7�!;�Hi9�g��i�t�9/���:�0�Y�N�%��dy��rnlu�Bs��o����~�CXq��(�"��@�q��#j4t4��'��چ7�&$��ՈU:"�\&w���}���С܆�=N$l䜣�px�d�)�L]����W���F����ފ��P�D��������O�	���U��@"�>O�J�zL���v�KP�へ�� "�����}Y~f����g��U���G')���g�N]���E�M�\�"͵��c�G�CZk�"�_�B-��IJ�Z�0���G�<�"P���?��8Fi>z�K^�b�ˎ�����$(�2#��v�qlkt��_sy;V�-��Ɯ, �Ǌ�,���?�Uَ֋��w��;�,�Q����7�uQ�	�������iM���˓m;Q]؉S��*�ˣ��~������h%���"ʳ��5�C�V�Lv>�{.�P�#����I�0�[;:��Y�w�H�b�ch�ZeN�\�D&��Ip�ì ��4qh��I�G40�_�D�'*G�d��r��K ��S�]�T����d�� ������Y"���5�.>Vr�م��u���pN��j>2�"��ʷ8����-ذ�V�1���Bw��(�rN��Ok����d�[��� ��f�gSr۰Bw�Wo=Lg�
1���X�eP� a�=���a����!{����K��Hq��@P�-�c�YI�0�R���/�N��dG��HՊ�kcs�C���j!�V��H�-�v�?�?�5���e��8��e9���k�������AE&���1���74 6>�q4��8P�5��Ϡ#\�b��Zz-~v�#��� ��Ԫ�x�w0+V�O��u��@b����:��^���f���H�AUԈ�n�����R�[���v�]m!	<|?i�ew���$���SG�i��n���:�s6-%F�Y����.���
��/�`�	�8l����*����>�g��l2IasB�p����9iƿ=���������)K�E�-��f����.��_�XgB�LeZ00�^�����n�cf�48Xr)���E���}ݚ�\��?L}u\T��5��� � �%RCIKw7J7�RR��#0 C7����tI�t�Π������9�9;�^k�=�L�Y�¿����V^V�����T�&�'�*�-��g�j�}G��0tr�_4�����?�gM� ��7�9�ρt�صڮ��w�>*;��I�p��Ac0�E�p��7��ɐ��i����o`��E #�ƥ+삾�u b+o�2�v�����i�(}��z!�`���n�V�))����A�cl��1b�!���;��[kVЁ@��
\_�t�s*��,� Xo�T�6�X���9o�U]�gt����[j�����l۩��F���h��^�b��x�����HӴ8���H�(,�f���(� 8�1q�UBO-�S�O9�g;��F�a+��-�4�VTy��b.A���{��j����Y �b����������U�	�0Ɓ�n�e��s�8��)��C�U�l~�SQf�XuWU���r]�����F�TO#aU����Uۿ%NӞ�5&b@e�����y�۲M�L5����yY��7�������6�z�7l��	�n��ۮ���q	�)�I="S�7�C�Z����˸C���K��bi���۱ܥp ٺ��Q�Ք�~�ϽA�����2���L�B��]WǛ�ؾ�955����|�_�HO��8���/ɱA2B�z�ed�c���m�[j9Q�X�ۀ(A��w� "�S�ۜ�5m��A�y�T�G;�L�M��8~Y|Xn2h5՟���߫�8�nr�2�V~F�� tt7yt��讎�y�sc�>0!sa��f8�G���[͂A{�!�N��v͢��Ϣ_͈3��'@��a�`м�SR��/�[���=� #x�h��}�``��Q����<^��H��C��
C�*ejDE�Js����0�-��Kv�����^̃T���K��Ş�Aw�]�]�hR��]�R;C�v��c�赳�����V)�)-5��:v����e�r ���-@U���@z,�ic<��p|�ʿx7��utX���(�S���Ӥ��L�������&̍�(u��"�c�&13������J��˫E�˫��ur �O��������L��PR-��Qx>�N�����ڃǙ��;�ʙ�p�ʕ��l�Sy4Tqq���UV	(6U��+G�j����%L�+��K����m�x�,���)p�*�qw�;	��v+D(�i�/�H$o���a�£����[�����!ȭO#J�gNG;R�:�G���Mu70��}�0��� A����y��=��6n�|�0/fTIv�qtt]H��<?{����;J��k��qh�ڣp<��k�s;���j��i8�R�Vc�TۥD�l2�9�R�yؚ����B�:~d&}�K@���$P����d��?�D�m`��)�SRkJ��(��K�G.r+B&��U��vKkkϬ1�}2�S�l���؄qr�A8]�U�MX��6�3r��^TC#�K�@�;�!w��JF�զR�N�7�_��摜h�e��2���b�
!yw~|��!;��s��F��N9�O����!j
,)A�3�L  �DDŖ)7�M���#"�ꛍ]}$��6ͳ����3$��zSTa>���1e]� ��ɳ�����E�"��9�� \%ȱ#���|���.O�k~ވ͗��3O�H޾�2���р���d� dn;��q ���R!�;�sjW�`�X!��cm�"eo$9�O��Q�{�[4����ԣk����� o������#���G�d�~���~;
&C��Y<�!�����&�m"���&�@b�k��X�����	��A��^0����g+���]�7^̙C�o���P���)�n����[
���V�s����f��:��{1�����~�l��:%N����f�F���FڣYM�!�{g(����hg1DT�'1]��'�c0	ᦖ5a崻��gD����i����d'niU�5��Z�(�o�!�X�|ac�7rJq�������w>E"��g�,��Z\/tb6i��� r�k�H�Nn���B�{��X�&)1Ͽ�0 ןN콩�oT�����>����q�0�d����hO��fxM"
Gb��$�����ʲ�>ql��_�8����%���sF^�d�߂ET�?:~]1��:�k��.������z�٨��c�Sr*4����L�-ݨ0Hw5P|��VY�
&B�bv!$���6�(���٦��?�J���XU۽ڞ�/�Vh�E����ǪGA^�2&�$3������R�""5���p�ւ[�M�����3�X�i���s�" �a'�G���a,.�!g��u�<�b�9�^�U5�kLa�<@�`+�n(�)�*�!���?�;9������p����p��	m2�1D1@j��`���F�	I�n���<��/�y�H{�U�6:���FD�x��6Kl�n�?��Zi�z=��t_�\��!x���~1"��>�,|*�x4�68	��� ��� �3�J� x��^|���g=շ�d������g�͂�@�f��N�� ��X|��\���" ����;�Ly��}����-zl<5,�pH���f=v��Pm�_�wuf���$��S�7pD4��"{K���I��.YV-�s|��߱#�iW�#��Y$��~��>�{��I*b+��AѲZ6���2�]�f�[��X�;�y7l��x1ŧ�\�������	ȕ[��O'f��y28SE_�ˌ?xBDr�y�m'�K�=��oe�i�|eJPZ��9>��B���T���O}�����X�&E��(�M����J#�wG�AL����]��!�g �y~_��[}�oa���x�6so2@<2_@�� 	r�=��~|"b~�����ҩ̌N��k:@�!��kf��f�i���t}�Q�A�(���h����u�b!�o_.�5Tm�X��\�Q!~Ws=�g�v�fGզ���̢�6���Nfs�� �I0���̻�4��?O��XRG��2O��gU�u�QRYћ�-�ן5*����efv��c���:x��p�i�1#�i]���g���N�����jJ|��:W��e�M��9~U�ED���dHvm�I��+�X�E�J 
5��3
f��J4�����^	�J�-��%��� z���k�~��:�eo�9z@)`����������U�������b��%�*ULgV�F���B�g�@m��(f��@����~���a �i+���~�{%��c�O�`��){�����A�L��G�خ6aΊ�������z�Ӗ*��G�H�� �8���7���4�8ſ3�>�0�%��j�]�8�N�[rȮD�G�1����\��S�{�V�+s�L��TwŨ0 �3*;/,~q� �d�p�3�s�������:~�b�mAf������[	�Z!"�J^�(�Z�4���C��abz��?��*Z+*��C���LV��X<*�AL] �H������H��Ub�.�wBhj0k�̏���N�heC_�q��n-��F�;�N��e���c��ƗKz��Kq�`����o�eQh�ӡ!�[������l�l��
�c�����<���6�^��I��l�1��u>Cm\ֈ����~�(%$��5q)� �+[#f{J65�h���Ds�|�וV���B�b��@�P?�Z�_~�_ ݗH��l\��!�/#O��˝�5���s�ۍ�Z�ˁ��l��#ݾ��E&q�.�U�����2D:��ԗ4�EN,�Ê��	��� �u��P8�j!�Q8�Q��) ��4E,O��NQ��n��[Ъ�!R� �|*��^q������ز θ�ԅX���(���s���'Dl���I�2�"�Q��e:zy��>.V�l~��s]ca㒳v{��٠]�$�=ڂ�̙:�%T���l�0����^��wH/]�\he�5��\Ij�����y�����d����m?1���.Z�^6Vz#U,��S��ߨ��5t�|3������myq�ZZ$\f̑��qf���K��r+ͦ����Ѽ	_2���}�����۝�,5G�2.�/AtqwF�t�R�\k�QY�����EHPI;D���IS�Y��u{w���}D�eCkN�])kyTz�[s"�E�J[J��&��j�_���E���i�+@T��;����0_�d*s�E�f�)>nr+��v=*����A
�VtK[T��v���pe7�}k$�.C}ʜe ��( ��/)��0{9����� 0^�d�z��&�>{�"#>�я8�=Pm|-��+f�t��M�ל*�Ǌ��N�'�=���&�V�0l�A����en0`pZ (o�r�K���������?ij��XPN-V�J-
0�4ٿG�v	�q���SQX�P��.��J�.HPpų0vpP����(4�/L�h����vu��.2N5p�uv����]�q�o�@ *1*~}����X�ru�n��ѭ<C��@Aa�o� Qw^�������/���[�Y��G_��X�[�[7�y��(��NS|OϺ辴�"$\�B�&�`5�m��/7w=\�4r��1��X.��?E�*��5�k�?zq
1B0����ӱ3���{~�邙?# P�!Z��J�x9)�$�������G�e�:����j+#Q�j<8����W��6����\K������CC��Q "�Sİۑ��B|�Ύ(�[��C�e�F^,\g,G}�B
���^.��-�9-������G��	ng�Z<u��ܭ�F�y�������� l |��܏��yGf�f;q��G�ctL$?$��%�������Q�^�%��Z�U�r �|�$8xL8����ƨ�S���ye�����(F�wJ�)Y]bP�C��0�(:�e�b�h����'�:�
��|�O��_G�FI_�֕�W�� 8��T��ۜ���}ۄx�s��͜���M�`v�;���E@y;W�ځ-Kb9�Ap�o(b�����aOL�y������3����_{�[���Ց E]���$��d<M4:/��"mj8b��|�l^�w2����j���մS�s#���pv�[0j���ń�}	����k�%���Ʃ����<u�i�?~�t(�� ;���| Cl���RRf��(c%�V�|ķ[�53���k�N� ��q�e/k�$6��N�d��s:d�]a2v Y���8_�8O���GO]X?�� �Oޟ���.0������~RCnnB��׭�Ɂl+������h��T��;R�xŏ�b펠H���;�&��,�eK�m��g�3�Lj�Kh Q�h;R3N�	��E�8|��El�IP�jh�'@��������9>b�<D�KbW;��Ky b��;��U�9�w���(����y�&o5W���<��e0_�,F�-�
������{�`�3=(D{�����:1�6��NP��\��r�����3pX{�T��u�o��g�+��I'&��ۜ�qZ���;��MV��Ԣ�Mx��uT�N�VSN���ԨB��.sV���\#�S�I�ҠhK��1,�B�Bg��V�Se��!u�Ľ��}v��u5Fl�gui#qA[��Cg����DNԔ������c�����oo��>}�՛۪�3�p��0����-z�J<`-�"�ݠ�ܿ���1��O�2�AO��t
Ũ���?"��acX�����u�׬�=ۧq��keh|���p���M�_�2	=AL,�q�b��2�Q̯X猶\;�u�jݿN��W92�^���@}T�%�K���6����&+=@1h��5�)\�Ӓ|CK����U%�ٶ���6�y�&���o�ϕlҲl+k�������߾���$A�j����t�Uu�J��LܮnK���'vDH�7<�	�Z� )Y�y!����O���F����e�ZQ:b}�/_�ZZ�_��Ȟ�SPZ{HH�j/�e�3��B�" ������gU]x���wջ���.��?�1�%�!��� V�E���W̦�~I�L$=H'��}�c�'�^��e/�ܙ���k�(��*��'��V��}�bBA�C�=G���o	G3]�V.���+�f�Uژ��8^UĊ"�����@�o�(�g
p������u��ZG�t٥���c?uA,�f��hgǙ�[P�?)������������=4������oFx��\�4ʂ�{oc Rc��.�;ڑZ���Z� �0[�4���X*֥���5;�;~�"�j��g�l�9�^R�4 �����q��3�v���s�Ζ��^�d:�'�Q���A-���)�Y5�j��s�/���I ��׎���4�`��gg\��X�xe��1'����A!-7�;��T[������?oz��@�.hg��[�����Ji@ɗ��x��D�
��p^��zʌ����ᥚ4K����4���럏���Z��Qѕ�(}3�\'�z����#o�Ot�U���� m�~2��#>d�b��$�L���+�-�F�~y�s�B���B�����3��҂Rlu�ޥ��'��>�5�	m�\�7
/
 7wՓa�E��_�R��ߗo�(<i�bU�ܡ�m�T�I���uNۓ&�Ŋ��l��o1�Շ}.�Pp~'�H���zz����b܂�(�zf
&h�K�j�!Ӣ�E�,3H��a�J�� �����5��g8���2C�=���&r�j�$J����̑.[��v�.�7222DGKO��5��{���DBTC�5���q�2{�h;Vi&�я�8ͱ4�~�*4��7\�n���f�@��Ց�ݿ���+��a9N�bu��WVW
����o��A�O��:B�a*���޽�aX��	]��UfK+��fS�2�:��Yq��'��"��O>@��~�p��<���R�*�/QZZb7<�k���-#�Ό��䖘�1��gAuufPT��F5���Fɶ�����V�[�����Q�j�n�׹�\�'ԝ��)��8�57��x��|c{�"�=�����kr_;��\1���PNB&�����:�t�w�Ȝ�	�UAJ��8b��=[��C������� vU�r2�ܿ;���D��P�3���<��*HE;ǎ�%&�f�c�h�w�X~���O&��-����c��v�jn� �l`�>xj'�+I��/�S�1��X��
�?�5F���}���U����c)|o�_�(�A����ZS>w�(o9�۠�]z���B���%@�Y�澠Nir��+�jF�}�G�1�R�鴂~�?��?�����4��#��嵰#��=���2���>���:�nHj�Sp�g?e��Ja��28,]E#_���y���tz|D���Y��/朊=��t���tR�4g����2��m����/w�W�R�>1v*h�h��&�k�����g�����^S��)P�f�ZHhsc,��ʖ͘�������	���F	���l'�66��eW �0A�ЗFZp�wb�T�����5��4�?\�-#��.���Ym���C��j���J�4������pZPT����0'�3~0�M�(�O�u��J>>Dr,�؀�]��[ �,�h G=���U��~��\G�E��^�\r�$N���T���C,�+�W�a޺��Ei1�W�K�&��g�Ǿ���#k_����k���+���Yvqѷ��Í�!�\w7�+��-�-h}��^���Ev8}�Ǻ�pfTѸt�x&�|�N��!���U��\x�cm��	>��垭�f�C�T'&.1�Rx4`8�3,�!QP(�Zf�"#Ɇ�[Zb�O `���g-���~���w�~S�A}�u���<�z#,��/ �����x�j�1�C����h�ܒL<��$�s�ݠoq�Z��e��~z�����xT���/�R7�da/e�g�5�\���$��1��o��V�;�E'�j�2̅IC���b��'�H�ZJ���
qt'���ͯ0D��^>��>c�M�n�����~.�%�9��\��B���Tm�U�h�t|����7y�h�Q\([*�ėg���&j�)g=��^���#j�Չ|�ڎ�EK��HB�4��;�{�Ebh�lyRj������ڛ����?,�*�\�AT�T4 Vnَ/Q�]��5R�#������o?{���0��jD>�����R��2��0��	��I�`���DKF9��1�D�N���k��$Ό�s6�oB߶�hW���2��((�*��$��mN�>��x��!j�W��YS��M�S�-ٲUdXy_��O��5ϦB�SFD�__�f�!ɫ~��,r�.�V�@����`;��(�8����({ N�nO��_�
<;�}�%\�gQ�}��J��?kډ"V���3L�(���PQ{�Q�P� ��K�:������bR3'a&���ߓ@���Tί��Zj��G�Tڃ������v��n}��k�?>s(��r�s��# ���@z��MH�I�d�Dꔌ̧;;k��u�7����d�����R6�j��}�U�O�׶[���{ETړ�^f�i�ث���>C���R}�M�^�g��!(T�*��{���^��������*Z��
���?�ۅx��i���|��+�۠b��$�9-�I�6 �7u��&z�m���e ���8��h����=O ��)cg��x`��.CB�2ڿPOm���?ў5����9�vrNo��W�-�^kr�>�����ؖ��-ݖ9{j̬����k��~X�3�nm&X����.__�O�7���+C�͛�5��<�.? ^�O�\e�O\<��%�:�߳�+�V�W�/|��%�9{�T]�IOO�ʜ��^�Wu�{�E��{�O�s�}���{?�@�E���s�ߨ'P�z��)"+��cBa1j� ���[7�JJ��H
~��yn��?�aD�B�~�%S�6��8�N~�?��ډ����r~��UO0[8$�g�G5\Ե�`s!�]%ך���.�H��κ3�HH]�^,2�n�ZU�AW\q@[�_Iۏy@��4w:�~^Svs\�L�.�-a���U-�8��wR�����1����ԚO����u����l�@�K��u��� �j�Y��쫁�NM8�ܳ:��u�ˈVA��l���s5����l�c?�т@��R+\�aȽ���)R`����A�`r?S����y��bą�ͦ,��ҫ�1�+r���ʔm��.+�� ��U�u�SG��p�J8��!Iv�����	s�g�O�u�cS��ol����*���@_�U�ۉ���e:�|��Ǆ􄷨�h������I�1���Ns�N�I�6E^U�Li�$�)X�9v)��Ȳ�oŌ��>����D��O<�[p�*/Zu��`?�%DN$���-�oLWq �)_cͩ����� x~��3oP���P����}��IZq�֥���h�����~qY�E��o�f'F5�o�v5y�979rlKv���]6i�`�b0�y��`��u�D�$�d.R5?̞�v�,���������n��'�c��AC�h��p��]M�pޞ`�5���̶�e���w�K���Ť����A�k}��@���E��N��c�ƭ�?�Ďl� ��A�0TJ��'�s/&�����C�jPv��'��Att6l���L˗���Z�И�qn��o���a�N�<h7.5UlƕI�.�Y\0���`��G��U�K/��9����K*�:�%.��R��-�[YoI�8>�Y�qǚ�?��;S\��us|��7'�oM���7
�\䁽NYo�찗E��^~�����w��MmS�R�,**%�v���c�hg�q���z����pW�;������2uУIQCrѣ�2q�2:T�?�]��v�Wdi˵�e&n�po�Uy�2�[0���uu���&�H���Z���ڷ�KÞ�ӡ���e�ٰ����I�kk�/���z��i��hk�49`�����A�����'��<�w�aw�;��t=�g�n6�+��,����G��[����u��l��d���ҧ�d6��!��������3꼍��>?��Ɣ@�j�NyN��r�I�p�Z�uK�)5^���>�:N*}f�ޔ+��jԠЧ���+�p������?�$��1J���l�aP�	����P�ד�a46j�&��� �1<s�REBx����Qt��D*�v�	�_���� *����rN�"�����t�����L��:��i܅����LwL�6���c�.�R'sZ�~�v�}�a�	��ޛ��+���d~�ȓ²������}$�v��V�%	��>OH�cf�|���o�@Y�?�9�{�i��6b��I��K�bw!�Â�Tz���86Q��Ds,�l�0�#����j3ԭ��p��'.MNE~�}ݝzu��O7M@��|�� �}T�M�.��Jt!���`�;,�!ț�O_�@��T<0�R/�P�/*���qϒd��~�c���?#J�6:���{p'_����m���tw0x+Ȟ��H�H��GvTC�t)pG��Y��c=�PN����EX΃_n3tU��q�B�JC���.��=�����eD�9�Gɔ>��T�F�D9L���|�ȡ���6.8�.L���,'��+�0?Л�m��"�G�폺�2��#�MDI�:N�f���i��oz'�|�B� �K�;y����F}2�Oo��}��X�X 0UCK$�����P�7��<��/>����G@�$5�7b����Ɖ�5�)�A�#O>O
74��y��E�M>Qw&��\��㬢�&g	����&O©h-���Ȼ[3��3�xF��	���d�S�͖���$�o�c��\6o$�LlX���^��&o1��?B�2��Zj*J��J�]�F�]h�j�����ש�I���u7��Dco�+�٫�Bo��Qw"�,X��R����æ�,K�h@@��-_cV"u�l�~?�s&�
����F��}��N$6_��c���E��ʍz��5E0�����ّQ���1j��-�&̭�G"�U��$�+#��w{J�?}=��o'�k{�c�+h��H���wV�C	��)�� �5'C����󳾸�&����kv��"K���/y4xΰF�C.F�G8���~����s.o�t�Q����<� ���x�)�f��6�@� ���QE�>h��@� t�����_z��I�L s�1�鸓��5IK�Mt�T�Q���� ocFz���]�i��䑶A �� D.�Y'C wQ�sg�\�J=3�T�$Wwe�t�"�7t���oڐ[A\����&K���++<#�Хs2)�r"h|ݡ�O��C����~[����ꮄR�A�p�PZ�P�\�'�r�:2�zw��<N����9P�S�֌�[ܿ_���D9}S�O�Ҏ+�[�X�6@���� �Y���WC�s�+�\�{':�W�N�e����2~�.��qz ZC6�A"�]�k��!���v$�5�7X��9� ;Ocg.ܲ��9��VC �}gp��B��{��ΐ��Z� |�=��oW}����?�V�拏u�e�W���� �p��bZK��hg�uR@����f��4���-�C���;Yb�~zE?!�R|������>!�0�-?(N���01������.�=��V��ƺ�R�<�E�偺�xx�T���#mm  )�Š���PE{���6�^��~�0��
������N����d�3���D�[X�!B�< ��߻9pՔe��X��N�M��������'�tW������[η(�)���=�|7�`j(�i4�-���cX�����.;	���O�ӫe���8�-%b7�͞_�$�vt�ּH_��5���Q]�����?�FP���9�e�m>%����Q�����h��1 �!x+�s"�����ط�?#i���L��r0��
~����H�s'�R���I]�g�N�5e��D�k��$ $/���Uw��M _5Ϙx�N�M�����\�fMK1GH���l�Y�����S���p����e_0c�����Z2RM�FR��򲃃���^ W9�u��/��n�8,R�q�q
s���E�Y;���oJ�:�t�a,��9���PL�Cm��5_Y�1�lx�u�r尽��1�)��6s#���'J�A�iU��u_���ꂍ|�����nyŦ��C�4 �ݿ���,���rQ������������#m6�G�F}I^}x�.8c�����*e��-�T �TM��si+P�!Xx:�	cn.�:L�ﮍ�'w��J7��+���c��v����%@"];�A��Y(ڭ��_q1U��l�(�NB��6��^cX�=dp6���L�N"��E�7U�4��*.��<i__�x�x����t2�~�"A���]�6�,�ל
"�������4d����]�0F~`d`�
�Y��Oİ�X4�_�W��M~�;;�}�o��-_�\�P^o����a�YșN��٘�����$E�&��S�7K��`J�W�=��}��O������$g��i^/OH�z {��A��ĵ�ʟ�?;jrM� wɕ��]OR@��t�4�Nl���֡���� �4��l�� &��QQ#z�W�6ܢm��h�?
�+�?��
4�B@&���N4~d��"�����r�r�MF��5G�X�'��M�[�h8	Sd� ��|��y2��`������4]g~C�;l'u�Lb��/vT�����'3�Úx���J�hF��J�U� 2q�S�3�<���L`�gHR�w�A��,>�:܎�.�t�������Z
����IO�H�]�g��F�j|q Ѵ&����@�����ߙ 'F��6`J͜ ��4��� �Q�H�1P�\rԠ;kb�;_Y��y�W��F�o?�h츜��T���Y�����ˣ@��f�<�5���11��Ps��`�΀��"�,!?�g)}2���X[���xpX�1�AL[�R��=��?@kQ��m�)�O��̶��O>F�'���k.a��ֿV�4��B���yJ�v���W��SF�"���K��*&n��P~�K$��]_2Nl���f�/-{�uE�8�ǥ��1��k�rAB%�mP`�DH ��'�y��y��?N3�E��{;�pv��	�_�� d��/�t��I����<�1��g�^��Q�+�2�b4�$r	��m�9c�[��b0yjȩe����14�A�	rXB��RU��E���:�Z$R��1�����G�۹�q �G"8
��#���B50�r(�C��0�E�TT<���$�j���fM��ɮ�y ��sR(�|�8��JA!�L-�	�9�(��K����I�b�T =�� y{'S����'�c����<��\��{?n�$�+HT�lNTM�I6��qV�5ۤKc�������<"�lLU�9���+�W�[!���t�@�Κ������$�@P�M�#?Qt~7y[����H��k�~��ޜrP�
��"]����������併��}������LoǣL���׶�JQ��)�[MF��cz��/Q�:��F�_Aw��{��wK� ǄO%G��!�'��,�ڨ���9A�c��3��1s���ihA����o��M�e]��7(��ˆ�h�[���䑡���"q��@��@B���^��N�]0��f��iҡ;�����?咶hّ�����5
)x4�YA���J|�_C�{�N�]%��rਗ਼�v�K��JO���C,Z)qNc���89�T�Q9/�����.�7�0*��'l��Vi���B�x�%��@�#�����z�qO6�-v��ʬ�<���y_ZS,w=��Z0��m�!=0����sG���'/Ɛ�E��Q��C�3�F�ssz'G;Hqs�s��2�y�U%�.Mv�PJK�d��ݭ�
���^kƮ�f6�&yD[�:1������s�㡒�յ��ŚM��T�Э�tAb��瘌G�����m�Uz�?�0�K���3s<�g���q�$�ֿ�3�n�Eoqԯ��5R��3�j!����Nn�]\rQ����Q��n��#�� �2\#�z�œ:��F����q���i��i�~�a'�*�&�@�	�c)+@Ĥ�Qݛܮopĕ� RC�P'�??�J8p�<��N���F1QL�tЁ4By����KI^�T��{�Jg���Yak��"���ۏo\Fߙ���^�����	.S�E���(����aEϱ�Jc.6a�_-��8~�ûT7���qa"��Գ!�cA�� "7F����k������ �$J-Nr���dҩ��-� 2/l�p���]��j�N#O���[)Q��q7��O��b7r���#��,;�����c��B��̧;r/K�5�h�Z���Ԓ9I���ef�1���|I�D�h��Ӳq�\�7�;s}8٤J�*dߚ݀�>�v�촭>�v�g 6/X�`]C���oL�{aT<gxiP?N�@m���;�72�<,�(b�6�-��(��r,a䝴�N}�$�g  �1P��T���R��`�Bl0L2���/ʏj�%�%��������޸����?w��=�x���e�ܟ�v�4E�aj��b�[3��Gܚ�#cu������>��|��h��N}���9���y�R��H��V��l-:Txc�*��M3�q-t~`	*-b��}mN2�ЕQ�l�"'��Z�����)��(�^m�_:x�}��åEE�r	�p�/����;���� �֮ߏkG �� �3	��e�G�{�_$p���=l�]��m�>Y_c��˪���`5$Qv�
绎�R5{_'W����w������5T�Y�����0��ⱞ{3B	v���d4!�;V��'#W`|��M��v,�R�zX�<p��6M�7w�|�m&sz5��1�q�h�LT�m��s'�\����w��K���D�:�n�F�v3#�4�+�@M�Z�ܚ/�j��{(=�j<����}�����{+=�������ӣ��sԱ�ML&�O!�Ov�sNи���h7�h_Z���4��F(�V�I�������:{�(2�Ip�~���%��ze�ԡuq��b����c��r�&���FFn���<�_x�c�3�o��b�ʕeZt�Ɖ��QAG���"��R'�D���uep!�)n��8���1@���kT���(��?�?4ЗH���t��=7�]�FJ�X�)3����k��򞓄l����U�u���~|"�=�[Բ*�6,\����W.N�Q/�\�11��� P��{BXZ*=qS�z+������,�
��ZP�v����z�^�7���b�.�����8�R,���I��o�d=,�A_[}�m��>tpȶt����ɜ���)���/��s��<ٽVӈ��i<'���ViN9���#�rx����<���]����B��(�ҩ�KM�
�����_zh��h��/�@:7P��o�с�e����4�M��i��ā}��H�m��q�so'۷���P�Q�&'�!�Q09��N��G��#u�
����:��\���������C-��ޘ#�c܀ț���z<7 q!�1��Ҝi8��i��f<ƛ�l�I�$v\�m`�3y�Τv��V?P�'>˖�{����y�+��%�1�!^%AZ`��pIE���}�^'H�1������7�I��X�&�%�SS��v[ +�F���B^q��%��7�v�!wjq=k�봓��+|~��+1�����힒J{Xg-9u��8�$l�zk)���F��
���W�]�"�*��+*Xu'��Q+m�`�=q�E�5G(��p�g��9�gK�b'X�������3 ���b��O��.�{���V� {�Έ�C��Q��;��˔�Q
�H��:��@s��Ԉ"|�#�C0����PV)�"���M�N�Ej�E��u����!v�a9*�m3�|�s'g�1��p�U;�@���SB����o�<w����[���(���c�	�cnPw&<���~�� "M��� :�'��|�ה��"u'�NploN{*�z����J6�jw�A��n�)�4�S��4,�9���ɣ<���cNo��&�����!֡�����t�jC�6��^�cc�#l�{Hw��Go~�����q����8}(�F�gW�y����{wj1C|�(�A�B���^�~�+,F����>�!�	}�҃�=͘c�T�Hg�v��a��i�x;c��H�-)rݑq�{&�?%��Yh	�܎�Å,kX|f�&�ϭ���s.�A�R�Î�Ņ�N x�Y�'�u��,�mk�We��L~A������?�\_�z{\/�&D%xc�˸����/���� e?L'B�����4W\g'��$��1�n8>?cյu,!�E��G4�KZ�E�b��:�v�*���Y1�P�&�9.N��P�Yc@�-ЉL��w�(%n�E�Cz;5g%o���Tv]���݁��\j�	7�����HUٙN+��_��ٚ
 �+]7(>2��% M2Twz�V��N�pz�Q�c�.i1/_�y2��A��^[�u�ih1¸���,Y{5��$�|���%Wޗ!� =h�;��m�y��l����(W�՛7~2�/r�/�����l�~<� 2Q@an>EF`��@G��x��lo@:p?'%�����p�<Y7�A	���R��R<~��%Ÿe�="��;j�HA�V.oC�Y�*�"^Qr;,�&e�xY�|�bW�@4�2.� �n��ˉ�>j���z}S�WZ�c?�?j+��zS�:T�ъ&u��%�O�]1ۏ��#�nZ�Ϊܧ�D��6v��g-B揫�@��*8�6}X&	Di�kD ���3��u(���9����Q��u��F�C���7�5G��G�o<�k��8�����o'W��#'�.�m$e��1*�<WF����� �9���	�|��3��)1��Ձ/��x�ۡ�eI�dwX`bO.������$^]e�Ũ�3�[�������'�+Iwh�m��7����m���F$�؍<��w�J�l\��P 9�̣��%���1{Y1����Z��usI��ќ{�����gV�4sOMM�`��IÆw���(��3��΍&���\2%(������V�kZ/O�Ȭ?��9[ѻ �ۇ�+���y"4r�r�j��xl�6�����0��ņ��>aw��I,�Ԙ��ͤ���� ��k� �t�tI
��R� �� �K��!���R��%� �t7�t�����~�ץ��z�<3w̙����+�/�G�}�_�z��u���ߎA��]�-��J���ǖ�G�l�og�ד3{�ǏՓ�J�E�l����R��>�����x3W�ۺ���}F�hc��.#n$�p�^�[�&��}�9u�r3�H�4�5=�<b�s���I�W�s�N<�̠X�d��l�˔%�y�.�7�1�e�XWg׬��z�X2�X���ڭPQ�����I7u�5���W�+�?"f�~)c��'�|a�g�)&�lH=5'�	���ȟ9 ��a0=���r>��nx�觺F����r���<l�Vt�LS�l�\�Eߏ�������s�)b�bXL/.ל���碩������X��mq�Y�H�x���e<-�����������zV��zA�R8q��p�m\x8��oLL��+`�'omXU��L�!W"��w[�ͭ�R[Q/?;�<�=�
F�ό�d��*/�Ӝ��A�\���D��``�u�(����,y��%w��Q��u�?7:C8��ZIRp��	���FFD�|����r����7�����ވ� �����P���w��9sq���O�h��sG��e��V�!�R�%�#�P.o�t�_Niu��w��G�'�@E�C)���?��tu�LX�o���u�l&'x�HVj�C|eE�7�)�|��0�����H�w]2޴i�SDNm5�C��yB��/� �\?f��"���Tz$�"���Rgʹ�L������vC�ֿ��v�D��=;X�����c�%p.�g\lj�x�Z�g����b�#�I�R�)߇�V@|���L�MO�Pښ�S��h�H��s��u|�)q ۦ�k��Mؿ����|_�J�0���m�C��~�%�
8�f�;%|k["�	߮J܌Z\�𫃎������@��&�~��0#�����S ���kwg؛r8C���Ԯ�J���F��g6�%°�K���KϛZ!C�T�0��hf��Z��j|���O�V7C�w52@�\����{� �0���W���S�P��g�;�=�Ѷd:[���d�K��6hE8X���,��ܹQ	a<���>5���R�Ss��x� ̍ �빑Z>rBv4��q��߬���)�z~)���� �a���h9j���zش9��w�A>!}�����3 v�����Q��' �	U�����r�9Xa��P6u�y0�G��7U�����a��Ӈ3]d�������î�أa<޵2�\�QW�x(�sj�=pAOGIv�),�����a�~Q��i��a���I�=C+�ɕH��3��`�'��ޅ*��=��v�7�甼���7�/)���s/�(�S��-�$x����^M�����+o���ʊ�����S��TDo�r��)�☚��TݽpZ+���f�E�L,<�.��2 ��7ң�j���D:�q,�:b���#��|S�/x�M�v7��`;��-���gcւҮ�b	?�!g���@�/!���5J�в6|p��mט+%9�O��>�Y��=�嶎|� ��}o��˒����5Y�l�t�5�*;Gy�_��w[�8�p%��/��CW��Z ��}U��ҿ�B傴���ځx����D�)٤�n����Oт��A��nPo7X�缨����e[����.���Ļ2�4+RI���"��è�Dsޫ��2:˲���u���Q2(g>�H!�f�yu�s���������<DnăKG�³5���QCq����O��bQ5�L�i"�������3�U��o� k%�P8'ɫ�����'��E�!�<�!��Ѫ ԶKR�{s���O积���/XNmg"���VA��=��s�8�1�.B�$b�.Q��29%�{��G����5f���n7����%�k��.+��}�}�`�����9}���k6��K�jH�2 Jb�X����	BF� "�� ������q��b��L*�>Dy��/��k��?�Sz$cq���E5I��m/�s�	�3�](g�֔ֆ�P�73�N;�m'f�3Ԍ��y<b���{�����A�?�F�-1�(���%J��;�%���j���\'WR��=$�;�AIz,�f���a>4x����̤�e�c�2��ynT�����$�GF�5'"e�'o|�d������'~񔳄!��O��=���.�f:�Clz���U��Ywm�Pl�v*�� \�N�ҥԘ^yu�m'�F�Y` V}�����U�#Y�:~�lI}�к������#�#��:N���$n��Xh��;/�kjY8d��w<�~c�����o_�ts>�>��Λw�9)xDS��я�P�
�W�A���Є�p�"�I����V�CD�H$�����X�Z���z�lc�3?&H�����s�],>W	^��{��|\���DRO�98Rn�xW���2Ѳ��@�t߶g�U4/?V� ʐ|m'��b�A��gy�nĈU#�
gr\�v#�nt�<|�z8�ƛ��$��NS�F�����;�0�
8�᧯�Ya��h�GP+L���@�N��\="| h�[`��P�����E��鸆L��t���l�7�	[JW� xT���ir�\w�,��^��T|`���"�N��%�7�����ݒ�����]f��C-�B9�t�7䊗�t��L�S�V^*m������������.�ۡ+p���x�uC��2�jZ�|�ڞd��w{�"�Vڸ�S�]?�������&ܝ�5f���n���-`�s!˲���|��o�uf3��I�T��&x��'H8/O�d��8{̊��P��φ���'��u*R�k��D���9#��.� 	����g"R_�^��)��>p��(Z�'�j!���9�r�=kvq1�����$i�O�V�7+~��M�H�X�l���WV��O��}yY���ۘF#�<9�)�跾< �`l6Pֈ��)��.;Ji�'$��PY��0@�e|B�P{ϓ6z���P��`$�f��p�����*���������C�\r�wdb9X{c�R$��]�|�SpH�P�w���a�c�h*�#F��z?�,��U�%�8�2�,���Z�/F�v��W�!�$��O���-3����ۧ��p�#xSh�*#����w@�1�$E�K2�**��|�FF��1��5�nJ�lM����rFCi}8�B��!��*P�w4�I�k����U�`�yad6���B!sq ����b�������˨B��=���f��	v�+_i�G��j�I�&�e��0O�����l[��Y�١:�Q!�~�����Қ��#1Ԇ#*34�r�,��5�����`X)������3?�WJ����d$�@5��<�R�(��KO1]�}�gh�
C����V��䷽~��-���ʆ�)�4,A�d��4,ϻ�f'�����Ջ
�R���ȲL�!�����>�#Md}7�hd�X����D%�^�D_��{:�xR�p��Q��4��*�v��hxK!�tEg�#?����!�>��w�ʆz�K����8�F�����&}��B��}������ٝ@�y}{���˷�C�iO���Ҿ��>|i��ǃ�Ԗ�6���ެ��c���!9�ǥRt��p�ecaG��T�{��p" ?6##*���Z�硚r{�ގ�=wJ/O4A,�9�欫GT���}ĭaǃ�m9�<�O��*����A�-�lI��ȴ������ <n�xH�|̡�J�ПY���zD����������t���pdcʵ!�I�&���Q3Y��bg�^���@��F\�#]����g�P�+(*|(Qj�x;���p���"�+� ${�l��;��E;�§�9�-'m��Q�j�Ñ횁ǖ�^X���'*.�Ü8��u�n	��D?|_�<���K1���v��̓b�g��b����p�����w"�l��Q��T@����=���;(�E������(�Z��;��|���[�O���E޳N��70���n�b?QI�[���]֭Gq͇4�w@��a��UՠܯY�PףM�ć��+�.ǯ$:������R� � ���vP  ݂ �L��Z����(�[� ���{�Lb��<U���\�����ȟ����l�̍/�,N��02&�:d����z�]��C���(}�C�իbU�<�|���4]s�}����Vk;�]��#��
p�P
jA�{��aGě�=6b(�Z�в�����?j��l���"I4@�����> n	f�><��isIp�V�*�?�WЂb�����S|"J����)�j�n�j�2������G�g��UC���`�������z鿡��|o�(��u��Y�
 ^��C��!�J�� ����"-�d�����-eۗc���H$K6rƿL�'��q叓�M9��/��((��+�ؑ�P����-�K��Q�l�_:�#��_�X ~����M���^ʐ�΁�E�y�K��5���R�k�T9��fE��1��� "��C �0�W&���/�g���Ն�i��C�Ym��2 ;��4��se�����#��|�m� ������ľ�D�{���l��������Py[.�?-��c�G�G��֘��?��Qc����2'Wo��x��ܲZ������Sq Ֆ���y���H~����"N�P��2���`�Y�p�Igh��3FQ��u��pv��E�#���R�4��Tm��dA���}֭����F�k\Jw�s�J�}�c���=s��8!-\#	���s�ԉ����?��4@ �C�v<�n#�2�ɑ��wT>���7�cr\[B45#>���,ԪD*���**�e(�����e!�>�l���>cC�}l���q�Uß��m+���?��Kpr<P��X�Lj��B��L�2�J�n�x~�_8a-�x�37�L#�4۳= 6P�_�#y���w���/?4�	)q?PzS���>
RT�g�i������c��'I/౰�j_�^��~�Ė�CZ��+���C����-���b[�s!\�F�̸�b����r�K��⑭`�ѻ�<��D5˃a���4�P�˨��u���7�[؝�r��`��#�]DM���ȁ�8#�`��s2m&��-�4\s��:��=�Ž�W��j=���.��9 j��멹��g���������N� �ՠ�4��K�]��.�vT��^�\f����/ܐawh4Ƥ5P�)��8�j����:�t�կ�>	�?�c,)���,&�%<Rx�.��X��[
BV����/�p_'�

�8������I
+	il��2��9,�N�}��1ȱjRҜ��e���n�Tt.��<���t�v!���=���ߑC�^"�!҄?A77~L�$����)����3��Ѯ��'r���y�`�x-�vy�z\����栾�������@��/�܆�1m&�r�|��Ы�i��4pA�e�)V��!r��% 8)���qƂI~�zX
K��̋����
p��#n�_�U�~6X%�'���
�5�I�٪0�v�R��O]�U��ۄ� ���)̓����T���~�w*����0	�$�����2��=%���8�i����/
�XH@����,���!�FNy���N�M��R�D�߉a��\���͑u� �5�̑z|_Im�Y�X�Ź���)�K�p������A7�}9
�Q�|���W�����B)<p�Д�4��c	?��<}Ӈb��l��h�~o
I�V�]��-(�J�N�|be�g�ǐ.{�JbS��t������\��(_[�U���{��E��_��i��ǈ��\�	]ܑ��k{�"�8_�E��Z��N[g	�ew�!]\D���$+7z�so�Do�����⠹5QMgJ��ꆑ��\I�?U��πE��)��rY���r3ۙ�FSJ����洼&�	�Wd�Gx���@�}�\Տx[쐣I�p�uj�2k��c!	I|x������	r�ی��Ƅ�G�����#F�0�Y���+E!^dr��iXU��gG�9@�o\1� ����S�o�Af�����-�� Q+��e��En ��vR4p�cȟ�1�,�b��s�{~����r���/R�d ��բ���/�Lg��6o��aJ�1�\rvƯ�>Q]8v|�f�Q�xIT��f�!qy�T�D�#���i�s�Kߜh�&������$��G�1+I�cD�Ib#t\��v����% �I�~�E��;>(�l���������N~��?�*�5p�&Z�t�>'��i�Z ����{�9ldKz6c;�`+ċ<��� ]q��}�m��WV3���X�q�
#j%�߾���s���=J�8ɫ0�>
%�A:��U�]��k�Y��U�+~�j�I���~T�*����1R8,:�|\�>�]�?i|Ɨ��̲��l�g�}c�!�R7�����6GT�Q��V�Y$��B�;S�ۑ37����l�c:Ŏ��p6�u9�f�8��R�{�>{�4��&F��˄ܜ�U^:B���3)e�V�0�3��I"�;iU�:T�B�]z���$�mԄU����E?ɂ*Osl#��h�늣��@��z�KB�}'��ȵ쮃i�'Òl�9X��RLwf�y��|u��,����g�i��Hݸo1Sȧ����A;���]{x�'�
�C������7"�$T�y���1E�u��9��RV�jhޥ"�j��y�y�t�jQ��W_��f<��u7���7q�ȝ������#C:�T &V���'���l|є�s���j�{!߾�o����g��,�P�I���/���G��i�9u�"kӆ� �˕U�$g�2P���J���5�,D���|.����u����uq�C�����c��y��N�ށoX��+1KIb
ޏifj_3��#[���c���/��^|�>o�p^̵�e��u��t`o�#V=�D�].
���gg���q.��P�e[�Y�I'�N�1�!``�A2����Q�~$ZNQv�~֞tch���g���ۥX�����c�w�6�m $�dqBZ�����h3D��޽��_X��D�7�Z��Y�_����ɂ��cq������l�D�S؆�̠Β���0q߶�0j|�؁��$�Á��\(��O �ſ�E��D)�5�}ڌ1n4���ʠd[Mi4t=�!^H���b�%�hV���N��G�^� �-�M�~�ZR}�ء�E�|�Xh���!�wm��z{H�����C6�,i�j�a�!Y�-��=������,:��7�jhəv��ʱ|�l��K£o�-X"�mD�s�	�\P�S���F��m��?3�
"t��,��Iǘ��̾p�����&@~��ZD�0���]L��M��=���l��Y����P�"��AD�+���T8Z6��� R��u,�r>3����w؆�������26}h)�g�pHd��z}2��+�R*��p�Ȗ2Σ��1@$B�mBO!�&�rɻ�r�K�աҾ�����~��YȌ��>�C�o������2B��7�Ή��	R�<��pz�>�:5y%�$|G�4����*�;��`���!)���S(f?���P��m�)�s_i^��:��2�#Y7��D�}9G��|n����&b)���G[}.<�ġx}G��|�g���������j(�-��Yqڮ#蓬W����^^�LY�N.��ʆv��
�l\�B�&z<�G�Ds�Ԧ� 9�/�N�'�Gn�#���Y��JI�W.��a����z�l;R����Χ���@۰.m.l�Dn�u�3$r���O4V��VG?���ӈ,�[�gU\�8��^W�������p�d�|^��4D����Z���
�1��t�J��q�Y��7Јbb;��U}��z��!�Z���}t��h�\�x(���,~�q�<R�٪z^J�M�(���uu5�y���.X\p�˹Δ�z/��H����X8��k���x{�� �+�����{D�u�c��4���w���S�M���+��t�����G�}�Y���YY��茔zF�ҝi.�a/��U2�Ly�IZ���t�O���Ò�d��˔�Ƿ귏�"�e�=�±#�X��i�TM�s��&�M!�.��{���Bh�ɩAJ���b�W�#��r7.`Ʒ���ڀɫqBV6u4�$.9���~�C��E���;��J����<�*��;*���=�u��R��a)��x���-��|��( ����wJ���#�,&�BS���M k�d�|�2p{i/��=So�#�]ߖL�4�Ǡ/��}�{�8�x![Xa�wz�
vz.l�=��YjV�Ռ�?���E��8x~�!_!̅��p������U�C(/�{dY]����NV��H���P�oZ�eO�ӱe
7>�#���� �E㴜P/��ϓ�u�Jn�tM���u���S�?����=�n�LecM ���Q��>��ld��&��̈́}�=�Q���*��C����c�tE�0�,P���U玌?Z�����'�1�1p�^��JZ�W��e���M��4�TGxU�c��K&_�Z�L��0������)@x����
�E�-��3��r4�+���4ZA5�
,�տΈC�\
�����}b�{�b���w�(��Y�v�岺��Є㾳�Hy�R��#����i����"�S�3��c��M ������3����
��A�,�Q>S�5St���~�
T���_<����w�~�+�NзR�|�y�Y�<�j˧�K�����4i�Z�mqƣ�tAW .��^��p��z̅>�h���<L�Q�)Y������C�ݱ�ki��JG�a+6(T)�>���;��G�|�Lmֿ���!�YT��s\���ѳ|�e�O�\�UU�+���1&������S�#])��������K/����.c$r%��jօ^�]��d�-�S17��i��vf��Fv'ZP��<qj������/U��\jB��-vN�0G�
�&D�xD7;(���êp�x#�puR8M�0[ZV_�seQ�M�}�"���͏R@�M �i���Z�l������־՛Z��m�[(3�o���Od��J6!)Gg�ۇ�|����T$��;+��N�7��=cF��ФƸ-�,�6�H�d#:��q�3=���,����ݞ���VY����P��g뺉�1ZG>@� vP���9�"��b�J��솓	ŁrL�o��!�ܞ��k��e�#־ۚ�ʀV�Ջ�nˌLJ�v��i� $�w�U��Y�Q����d��lb�<�e��/ih!ĸ(�UP��}�j�Hx����`��#�*OMg����(��{B��=e|���!��F'�n�h��X�^X�L~a�%����8T�&5�<�:RQ'm-�|���,�^$�}��x�.J@񖥩G/�/��'�Q�E�2�%u3�QH�ꀤ�H@I���ض��C�V�eѿ	d2��_Aj���x5�P�sc�ݙ����O�\�B������'����\��?^�=Ѯ�����/1�����j��(��m�clZbˤX|SZ����e?<����ʆ����km���Z�I����@I���כ�#6<�U'��%��U���M�$P��3�����C�Zzx��HG�GXA�mK�d��9��t�h�c �Q����lt�U��8E�=�q�����J
������ ��h_7�&K�ks.����ר��w�@��J��(�h�.���lVX�C,����R�pe���$n��3y�Kđ�'�l�VYp�bT���"�h
3\�"�\��B�HƜXv���vB�Xn�+-�֑ncI��Ф�#�o]�Ur2�n���[��^#]�l殜�m�wa��ůJ�3A�f�q.Y�	����[��:�R�~.�_)>o0˶o��U�eS�X͑;�F������k�8���hA�g��k�m%�T��(i�(�z\��r-��^Ǒ�a�6��VN���߾��?q��v-a�C+^>�@�AjPHK���)T�8�3B�G��C���T	�c��"��mw�����F����[|�≳*�o��u��P��oy��@�A)iܺD���݊mk�7�S=2�d�rE�B�����k_Q�� j2����LtR����"������~G��X��V4"D�e;�y����4��4��K�Z�E����X���CÌ��1��v���_!�N�3�֚�"G��*��'���s&�F�jaI��F�O~臬�B��-���)/-�ۈ�B
� �J%��P��z�\�7X�^�Վ׼�_��N=�/�7!v
Qc�^����|'�}�<�յx�S7:A-���,Gr*U#�W��-����:��cw;���F�XK� ��H�ȩ��m[�K+N�q���}�#�C��27����6��͌R����?��7�TMV���4 ��a�9���kc�r�z�L�0�aT{ν��8�UY��e���8PH8�1P(��d`�iyM@�+��5r1��&�&�ݯp��"}q?R��� Ӊ��8�ƿ#a�\?⠣�*&4��	�2� �JG�r��j����;���I���>��ֲ�Z�X�
����I�t�~��n�
�Xb'�I`jH��[=�8��tCTɣU�Y�'��pp�wj&�s#�o)��y�Ó��p�#Ȝ�'+O���(]ޢKl�!0�"�d~	=|oe�R�75���p��i'?�������őh	A�j!�E��������2r����-���5q��/衫�3q��F�-K��`���6����eL�6�dafp�� ���da<�/�٫�s��Z�(Q�
%���Y�ɚAg4���hV=��%��6������sӹ,t�^��g�]�����;��R\�a�+,p^�����IA����Tß�Y.��8.�OJB��GJ<?��&HZ�5D `�=��&Y����N�G�N�F��h��;!8}�u�<+����3�Hb�-���p�n�7�rK�k>]�=Ω+Q����$�,�}�͞��j�2ॕK;b�#�MR���S��Ֆ�j-:�r�J�+��l; ;w�L/���������4�1��y�X;�1��T^� �����2$)�(ڶ�D��ma �j��:���^�^//��lI���~�19��04�����8C����{��[1j��"B��r����V�z�	�V�����C�=�����5��}��$j�j��!G*�J:��#�aۉ}���~��/�q���Z��P[�9��df�۔���%�(�&z����o�� ;�C*+�&g\�(i_�a�Դ)U���<4��J)����� C��8���q�p�YPcŚWɄq�:��R��n7�	{�K=YDw�ͨ��>��J7cu�_3��Sk�����y�3l��۴�f�1�r(}HܺL%
��0�:������$Ьt���YHF��lM���;�K����M��8���6��`��ON�o����~w%�+we={x�)џ���a
�<ip%�+U�dv����a��2.j��l��8b̐�z*Qw�E�D���!��_~�!�L����x���'���PG�����o�T���c��W��z[>B|�\����,g�1X�R��ߪ@?�9_���v�K����8X쮎*�+	�ڢ2l���s,��S����� <���)q�����Il��!kR�1B�]m��A5��豽�߉�G� �Bt�d��QN�Z�=��n}���8��I��6f.�����z'6�RM˔��@�!E@�4���>c�XX�C�Z��M!����q�uu
���l��&���HՁ�̈́��S�b%>F��Dҫ��)�[Y��0*�W`�_X� �4����\�7Z�C�G�m����;���|��;l�Eǰ�,� \�\_g�9�0O�V���������	4Ķq:`t<�����t/[���n���0�S	�) �H8+W����M��@�l����-87�Cl��,�|>x�e��:����h�C��ٸI��8�o���Sr�/O72�N ��%Z��Y�UM�Y�;�"=S��A��ąz0)�|~ZA�?=��e	�act���n7���;�8�󙟃ru����#�D %��?ꧪ�g����y;�¾�as�o4��)QزB�ps�I�au�VR�MC�7�]t�W���`������G��Sϰ��$Z�To��+v�:��e��&�C�q>D���p�U켂�	�ȣ�oG̟��Т%�}�L\�o``�C���vo:��>q����\����d��=1����U��o�ly����z�2��t�+�7��%Zrw/�|��ᠠH�{�Zަ!�'��IR�J��x�y�x)�P��J����"M�j�"c�@�b�����W���`�#-w�K�r�;�=��Ͽ0 9"�@GWh�;�9����U؛4��+6�?5c�WG~�<�Ռ�'���M�
�o�-�O}��l}���eFAb���"�I!#��_=��w7�ߕ_e�J���&#R-ȯ����d�P�xi���E��=ɕ�#	n���i�l�Q�BW���~?�Η9Z0�y>�{��v���󺜞������K�Xp��J"��C�@�����&@t]6��#	̊i�X�yC�48E����݄��h�n����?o(�,���]O���׼I��xCz���/�����׿�O~ �Q�Jޒ:k�i�<�D���L�|�P2���RW��v��țkC'��3�s�*}o*�~~���K�[g��y<�}X��;!���ŭ����n��3�>$�t����S�Bq�F��4Q*��X�U�od���@����W��Aċ>��(y����[b`���)�9�b���
[�V�J�
�]M"�:ET��Y���5�$ѻdr��Q���(��#�� ���5��@0��U�jIMV��E�:�E��Ws�	0	i�Ǿ��� ���S���L. �ib���h��?<d�P�
�?�y������x�;���_�+�:@]���������θz�2>�a��G���c��o�`k$�O�����);.��\�B��_؛�b��#8>e�ی����L~�^IoJ���4�0�>�RϠ���"�}�Rn/j��T������X�����D���1�^b��I�k�!�Ǖ�������*?;�*9�$	~���֜əUG�ڙ�O׆��Q��d�Q'� >�Pґ*=V�c�I2���}���HQ��*��Ux�3F5N/|�"��(��nc�ٚL'�8�����o�u��H�,c�����1�7C�D��3]�>|[�=�)�Z����"�[�vh���Ԍ͠l�T��$����\��.}�2L);�7K`u+Oz�K^H~�Gv�S(��1��ϧ��9<Z$� �2�^jn���i��p�ɩ�^�o�� ����	F�����u��؛ĵ���OZ�5�$O��&)��Y{�E=b���$9)[]�0�S*$��o���޼{��%~}E��5PR ��#{5m*�S���n ܼI畦���g$H|#�a��\0���/��_�D|S>p.7m��ᔤ 4�'[�8�Y����3��U��v�D/ɼ��cq��;�"���-�E}=.��F����ng�4�8�I@)�gh�=�r*;({�)ə~y�f��dhv��������ԋ�=�Lw�?��9uTy�>0����4zQ��1��P��*1W|�a���d[��{.+=�Ip�=zGׯ?^m�'���q�T�c�	�l��X)k�,k~e��l�l�H[�l�bc��t]��h��9�h!F)T���ە͔�Ǜm�6ƿ�"�T"��F�Q<�x��6|��U����Q^e�J��6�b��XMs�z����/_�z��=��*�I���X����=.����@F�P��J��=��YQQ4�OU"CS�t�S[��k�TG������E� ^�e�VBZ�LTϻ��+���͚+���Ë����DD�j���� Q�����K���
�5	K��Qְ�I��������o!�~X��Ԁ�14�'0���2�~�r%�7x��`c��Ȭ+�����\�K���L�<�����J��Q��p��(�k�J_J˗h�4����h�p���#䅬zX��V�㹱uS�s��mU���c1�YY�n#����yS����������*G�w��5���ݗаj\�H2�{�N��+��R�ya�J�r�q*X�	#�l�M��j}�a�d�U��S��[�w�*��Y	����oCDh���zoyU&�b1/����l�!�9�Ǹ�4g��)��f3�������OO5��+x�[�% �=�ѸbR)�֙w����S%/ƃ�څ8�xU�����_%P�|I5��g��?�|�W�⹭�;�k���$BN�O@�;��(q�����D�o��~�QzM�_�-�)��24t��]�`��m�_�흎5�V�Kg�J���2�Ci�xn\n�f�G�2��ʇ�D��_�F���J_�:fU�qm�f�2G��FeO������DHu���\*|f��g�ݻgt�Y=<�h���K���"�U�4<�ܮȽ��5Y
QJ����+k���1�ybh�9��qxe3W���Tr/?���J�x�[�␺i�MEm���j&E��`X�/l��S�Ä��;�V�1�����Ξн'�{��+?�j6���:�_��c�5�7����9Uʁ{���s9����T��Aƺ
>c'���jT��e�RCƦ����Y!Y��p���?7l��?��DI�����\���Z'���-�I�>�I�UnR�7\��5g�����d�=�sZj�R�7�W�#{�@�lׅ�p:�7�e�7��j�S��*v� ��F������y(�Dōz�gesɩ�����Q##$�n�钴TO�Ms�2li��>I+�9{�ED��~�-g�$S2�OS̤�
䍉��d��e�?�Z�A����	���}.g�2������X������o��s���U<k�8�'�q.������&~bv��ўc�'E��|��^b,<��0�ՠ�ޕ�׼ �2�!�#�4�v���3Hn��:.���^�p�h�(Z���ܷ��%`Kl�Z�s�O	���~�z�Z�M׎�p������S9� ZY�U���J>�C.�#zb$|	9��5��R?�l�
���]��	/�ٟ���`I6��^��r��<����mX@����B*4	��fQ��hs�C�D�f��Ww߾����Gg)i�au�<sr��*�;1���#�&$�
�6����?�������+�j�XIM5�x��<B^�CJa?[d[��ںF����^�-K��J�4�l�S����k�P�\�[��R����#�.&ƳV�Oú���Ui,�(Μ	���,f�#��ʀA	@�������;,5��CrAq�%�^����JWU��6�]��/}K�s���^��C��}�V�N�nI��k���f�d�X{�&>���_� 0�4��mX�Uϗ�~�J��nYĻ~���O��л���w�*4�e9�>g	4�?��H$��ym湧0v^�f���&-P�LY�\�췱�����&U�x�,��EJ�N�P������|����/39�
J��������s�x�q�C��hm:(���A��Sw���BuQ�y�D�LwL�O���UE*��}[�ż�E�p���b�V�G��m.�X3pܫ>�y>�%/Á$C�������W&S�����/ԝw���0]O������D�o_f:Ŏ��P�=^P����Q��o�Ȯ�Ѵ)rkkX��^�4 @� �F'j�>Wz�9h�����߶�該Q�캬�I[�=!�l�����_�ƮM8j�xL��Jՠ+_3���r�ܹ��-K�Y:q��(H����r��2�j���5?+�%G>��� d8��qI����-����"k�g���}C R�`�z����oƮ��_®�� j�[��w�+j|�n�@�d�Q��pLF��g�4DG�߶��犚��+�Q$jn��ؼ�,yMt��FX���N�jz�o#�H� e��ٶ����[V٧T$�ܱ+lU��?��A� �����ߎo?9���g�}!v�c\z�i���qq=��&�n�F����y�&]�v'�H�:�1-��Pi�9%�
�o���,֨(r�s�V+��{�~Js���/1�=U>�E�W��&?�9R�&|I�V�/֬��R� ;�/�hEYʋJ�~������j(b�*F�C�uKRk�b�/��s�qn������w׸P���d*<O�1m�_�$���b�
D����$���(
�����ˆ%��8��_���J�y���U=��+F��x5D�V���wi�?k�R)�Zq��y���������-ZNZ0����ܬ�h~AJ �'._b�;9�7��p�Mo�y	��#�rtū��:6������	�S�j�._�~�MkGP^��w������uEd�r(*0�B���)^L�BVP9�0��i��=�uz��)~�v�f�ZJy�`��L��}������!]t��U��5�	LR�o�Rh0�((��V����wF�?$<�2K w|�5��x��:$P�dZ��{1�0�im�dR�M�����p�0�1 7��WJK��o��*	i���j ]�k9}��}q�ֱf���M������%,յ�u�Z/������N�a�[��
��HŢ�3=�x��6�:�o�E&&I�����j�}���UϘK^v��kG��hn��m�Ӓ�h�X�8�;Q����߃/NEW7��)��i:��C�y�|���$Eq�L�WaOm�4jYT,� ���_����BX��Ң�[���`����<?(T�!��vOcĺ&��n$?���ְ~���PC�)ďE�?{$�~�KS^���_�=)�"��� ����������^����h�d��*kZ,b�s@bӃj���:(�����[�?C��܈�C�A�����v�:i8�3�@��!?{��︅�챻�1ä�x��_�&lK#���W_���=����������R2�R�ݩH7��R�C��HI����ЍH�t�����f-��0����O����7o�'{DJG뻰Ф�`xVVYȮ�?�	��W�����k��H��ϑ����k��N�(�;�a-6�H� ݜ��TT�Q9`xIdӊ�I`�RшH���@@(�N\�w�LK���:&�T�L�&�c�S��0���z	��<����[U)}�w����<U�y��Z�L�t���<lܛ��|h{J(�k]lp�}��V�;M��*�'@�e����ڀ�gM�gF�Ly�j!>I>�����V�����2�U`��r��e	�~�:�TX�{�U~W�`�հ�Z=4Ht�h%���*g��Ap����鄝�O{�}\�A^Pt�+"�凵*�f�v%�HW����j�y�� ��������K�y/%��ޅ�پ~8���fO���&��É�M��D�B0��k��h��qf�I^n����[����'�
�ж?y���5Uwx��������y[�H9|��Zwjp��H�]�����(Î���׫�i/�U.	��[��С�`U��y[ۖ7)hGn͝�Ue��S={2�)���K{���F�?r[W�����2�����YK���<V��x�>6\Iot�Mq9�yN]���ܰeB�/��$��Gp虄���0����+����4"[.8�*�V`�Z�B���Ք�е.a���|�)�a,)��:6Ф����]��C�w��e�OP�� f����{)쌳�bS�^4�R��ER�;Q�m�3N�#\���垞ܻ�7�Օ��3��D�_�����G��*��7�!�4�=���=���h}�a���Aj�o����Q<�GBeg�P$��J�2��0�P�?����m��K��:C������]}�m�C����e������u�?7z��h����<p��ݪp��l�F�}���1�}�g]�3
�'ɞ��wh+�p�0
B�衸5���N��H������:�%9�6O6iY~늪�R�,��D7���~]\ݟ����<������@;������&��vVt�R҈����S�T�n�<^{��A����ׅK��!��?��J�%M����6f�U@���Y�^{f�4Qg��@\����}���dg��"��qI�^$p��I�F�Ȏ߸^N�����悁>%7�o�+'��h����g���W���dE�����eݷ
�R��Ō',���w�@�.��\�	12��r!2�a�f�������)�ƒ�=��d84{T"�T��([�z8��5�L����Q���ګ��I�	R$����&���gӐbYM���������#��
�U�A"�/�q��&"�ݑ�Ί�f5CK��2�\V��	�
t���
,l��W��P.��4����6�T֪�GDKB�/h�I�A��D��w���;KWk�uJ�:�t�i�Y;�� ��6�S�#�Ǩ��NiH�sz�F���N���s�Gu��i{�u�@.L����UEx���u�6|���0.3�ԫiD��E��HR��W��,�K��ZP��[��L q�Z��T�l�L��oB�z��
R�" 2�2\'O�V�.��H��L��4�M~��L8�g%ET���
c��Z#�'��� ��p�v��9�oЃ�H�������z�}YjH#z�x��`ά�Xj;j/��Ϧ�Ҽհ�YBvT$���B�5$طV�T�Nտ+aԙdL8{��� #��?-\X!A}��ٰ��r��;��$w�	�L �;ۋ<=�t_Pn��֒u^@�������	~�R5��-?�p�C���7�v,б5mJ�7�J8����8Y�+�ܐ�#6��Եn�5�?���uҼ #��Zϯi6wk?�̥�� �3������֔N�w�$�h��k�36�����հ�: ~��fO��� ,(�}�<��w�mN���ԜA��,��� �ExG1q����P�^|���zDt�ly�R����h-���p�^�*B������C�(���
�UF*��[3���(�6���* ߩ{������)K��	Rh�C����� �}o�F������@����{��2�B^��z:k��Nn�3,��_��ʴ�^�h���*��N3��яt�rY�l��Hn�G��x���V	$`Wy�<_�EzT��]��Ԧs?0 �:�QOw�4,�i���r�0qȔ=A�%�y�p�(J9�r��,���I�d�+��l,��,��B����A�T.A�A��p�֦#O0�9n����x;zZ�_޼����!a�	͵g��oi�)�����+~�r�O�����YU�k�>��浩�C���7��7��W+�ޑ�a.�HA}
���s�0�V��%[�W�|hݲޚ�߸�NfFp����F�=��	t�&q9���f���	��}�e�1|�
.~hW�I����8��x`����-R��&'A�3$���ݬ�W��/�*��%����~�p-�\`�
꒿�}w��~���(�ڞ�lԂ�!)D �9�JE�o���b�0��!�w=�$e�ܞ���aP� �;�vnߗ�����.��j��}�5ݯ�C�Sg[� ~i-!0!%�{%|�Y�q�_�z����r�wCN�3v��n'�Ɲ��G	����Q�-���'A���\NnB6;ڴ�	O� i<@fн:��sPP�t�0'<'�j8x����':]7�s���٨�rKiH%� t�i�6�׏�;�r��A���"�(s�D�B�d��2D�Ѱ2}x,fH����0'�	��>��-D�&�i��������ɐrY��ϥ�ł��e��j�(��d��e� 	oᲣ��[�dg������Bݠ������d|Q0�p��C���Gp�����Jcn��нݯ&�{���ȼ�
�*;�Z�2ip���x�p ��J�����o��ܖMJ�OjEy.L؋[�Q�tg��KE>��y���9�mT_f��V�,Xm1EG
�����䛽/@�\����s�&�2մo��h���*��fr��;�C�!�x�酌�ĖahR���M_BY�MHѝУҒ$����d�
�/���n8�&�H��H�f��wJHx#��C$��t���k�(H�6�#�z���W��3�p��%d�@M-�Wٸ�
Q��v8�1n�ژ��8��v���3Slؐ����m�gR��{�I�G�����;��@�~�<i^E(c\��BS��v�\�)�;�:b�GW����LL���s�v[u�־��U.�pB����!PO�ϖ����(`���MΆ��)���Q=������D%�a�w�j�V�J�̋�p�S6�D2�-E_���*HE��{A9�`Is�	�����~���S�S؉_�sv�� �f�顭�G!YLpQ2_ٰ�N^��Hr�n1��[8�߅t��;eǔy�xo��	��.$�i���\ae�_���֗H���$_��~;N�,K�8l��S��y������&��ؙ����ggRٶM#��CD��F멾u���C��A-��7�Z���.��04��A
��r�6��	Yd�̌q��I���S����~PY��\��uƃ�缙�����72֩G}���QƂ>t�_�/xE�e����=�ρG�/�w���;�����DIU�+�/�k֜Ï�������a�\]�i T$/�B�����wࢄ\k�:�����{�޼����V�G��W%�q�y�;A�@Ho��Y�$[V<=+�Ok6��й�w���h���Bl�d?k�,x����"X1Lq���YL�*�\�X�Dpg��/~<�����TQ�Ζ�(�碢�3Q!�Ĺ���,C�~Wo	]���&�A(�٢��A��~Z��I��%�ݪJ�	{��A[�p�y�W1|�<����ҟ2�!Ð(�S�x�.��1��1Y��(�G�iO]�&�~���妀�������˟�`��Nj=��k1x��}/���L*���d(M�Վo��4�g�k�ZL�]k�����*kA��f���Mz�E��	��0���0�H͔�Ϧ�Q���Ad�a6���p�ZH��QﭺOQ>���0��~�OG�	��Ő���*6kl�76GpN:M|���Kh���Y������F�҄���Ӊ7��[gi��A3��ϐ�F���+k��eD�C˴i%!Y��j��eT1��������c�j����L�9,����������]C�w��ƫ2wK������5,a-y����S�qs|>��������i� Vy��`�<�����p,�fD�h/�g��Ղdw������o(��{����#^�"w�'�-l��U����&�[wM��]3�~�p�����<�K��8I"���a�t$��u����	��IH*�E:��y^���9�6n?|�&O`=�(_��e�/�y��_��x��5�`���l�7UA}͊��CQp�4c������Z,���7?�<2�&2Iy9�
������n���Acc�Ew�,�}حVo^o-�\�.d���۶� 	�v�G�raXc1u���T��F���^�Ԟ~s7�=��j31��Ǯ˞��wOە	���� ��,�h�]���*�3���+#���O�[�ܵ=d&�{�KP�=$ �ʕ|��k9X��W(a&�.����?ڕ]�=TB؏��'i����Y�>��, 6&��R��{Ԓo63�i�����las6���ʭ꾌ƟZG$�a�x�W(��o�be�Q��*o<O2�a�B�T$7�7�\���k�Utz�B0��Y��WcN���Ԋ�,\���'�<û��Q�Ƌ?9f��C�����,/Oy1��KskyI	�e�_7�j��Ek��5�^6�_�v�2�)��zV+o�t�M�o��ߟ���������I/}�h��|M��I�[d�f�Ŗ��{ѓ�Ajbk�3�1��n�"˥�r��u�@^�.���R�1��`g\��L�=?c�b
c�d@y���Q�M���FI��b�\ 	���%&Š���
�c�.҇��2�����.��f;R��e�����$�*��MLM�r�koz�Bg���~)Z���Z�5q�'t��7�>�9�z�W�4�H�fc@�,�bl�	�܊���Ak�-^LGY����� Qb)bE�TP���Š�Qh���a�n����D�ނP�z�-���i��s�~�<���}�;&d��Wf5˶�
X,�\��b݆��$�㣣�#%�u�:���b�8���7�ނ���?�P^�<`��;���f�G�&`�p�(v���&��&��apU�Z�g##M��ex<���=�&���b�G0+?�4�<B�^���i��[���	�Z.�o�1J�<�x��M��q�G�c��<�HBʻ q��	�G���^J��q���l�]W�_<���RK�������%Xy�h��%�A�}ٱ��׵���?������im�vN�+s�����c�Tꌐ%��Y�ρWR[�#�>n�w�>�^ɲ4y{ŏ��O�	dH������93�g��$�j���aC˫�W���ӂ�;��K�/���݊W�G��b��lI ^�X-�mL� �p��m��ͥa�ʓ���+aYq"�&�v�����@�.&ܳ�7�^��V�bӑ)7��?&��W���u�#���ؾ!$���4��
]HuKϯ�T�ZI������Jw�4�=eip�A���ɱV�I��0�4��S1v64�S1�|R���Qa�MG�ʶ�fɠ,G�FU��\��K���Nn�7���Y��u��j�/����2<�[AB��d/8t�Ύ�e�"ܸ�p�b}����q�~R��m �.SiL�+�=e\𧔤��;O�|�g��*R�eM\�Z{�����34����Ino����H(�-^�����e��ۇ�Bc�u@����������[�pRʅZ��>�=dG^�^��T1���De�-��1�;�Y�Ծ.�f�򗏋r�`�	2��.� k�ɜ�� N�Q8ʹٲQ�ޮ��ħz:�ܶY���UD ���`��,��:��u}�hP �3��&���u4�QA�zo�^���F���5�����O����u�=bV5�*�7��x�f��8���!M�*Լ�_��Z�.�*�F9ps��q��My���%Tq��퓖j�r�"��Y�ȴ��q��A;�쁉�T��A��G��FT�薼��Mzh��i?�����c7v��EV���K��y����(��,��,���R�I#�xE�ˮs٣2���=�eg� +�5�記�7�2��e�p�A3�8
�R��T>�늕� ]lY��jƱ�ˈ^̮5A�a�_A����Ƞ�@-���J���]G�w{�[�=nLtE��L](�}��Z2"���ݲ��h,({�-V��u{Xc�u $+K���G����a.���I��z���@DO:���j�+`gC��D~R�4���R1��8�%C\0e��㣕�Pel=���ΰ��ٍҩ��Y�����f��f�OzJ��bg�O]��T���T5"#�R~�բ�:Q]������I�6mƖd��P?�����^�
'r��&V�2_�ܡ���W��I�\s>= I}*�C��;U�]��Tf�;R������cZ1A�����[4�y�kκw/<xAv��"+�w�9~������!�sw(�˷e��O�8�ؙ��s���v���VV�����`����	�x����-�����)���|�3|D�'�����@�N$���-?j@�O�LnH�(Ś60wo�*�.s�]���`����<+�:6�w�S@#X���)ͣjq]�_Ҿ����a����m�T� ��v�ʄ�t�W�͊^����ʺ�m3�����Y���Ƌ�����>�g� �j89��ڢH_��U��)9��E���.f����#/$Q����p;Q�Ûf8�rQ�3J h�Q���	���dr���q߱�;���0d��J�*����}N�V����Dk��_�7I�/��jAl�N0���F\*x�R���=n���c���e�]0y���^muɄ�u�Sp�{U�gQ�����+�=��|xj��Z#յ���M��k���:=���z�Yd_��h�C�Uw���qQIW���<Y���d�&����{0�M	)��W"8�1����r\���I��{������ dZڏ���J���U���(��]Cs�<4qF/өi(n�5;�(�;����-ߴ����XRrǌf�Wn6��gP��vطfԎA l}�M��
�D3�au�ؗ�ԋ����d��p]���+ �	��,:O�
��Ļ���B��Cf�`~E�lIS��ؠ�>��t�e�Sl}(���JF��HpPvn��M��̕����Q�J���#��I4^��\��f1=����q�2^,b�����^Ѩ��O$�۶��]/m�*]הS`�t;[�s)[��ۭ���M8�ʿ-k^k��Ę��|�Ԧ�� �Y��nn�dF
Ȣ����pG�DN�0.�������5��c@��^��B0 Xr~z�^��
j��"�#�X5Aq���:��t!�aSa��iĎ�X��]1��S�U�Q1��|�'G��+k)H.��� ��V9��V'9	@@��R]\^Jo�$����W���v�������R�����?[��/�DW-;�� ����g�/������Ї[�<2N��N��v"��_�o�yC��6�o���TH�^χ��XdM���ˠ���S"�C����b��gx;M!	��A[���X�[H���bW�!��Wq~<��۲[�Q��'����nض���y�"��# Y����h�*�2'D)��3��MsBeW�"J�f�L5���X�L�ca��|أ��1m�> ��t���-���p�3�(��C��N�ȳ���ӁF��H�X �P�[�+Nƫ�#}��
'�P0�J�� ��`o�3������Vj���r��)���0�r�Sg7��\�&���iz�X�R��a]�+PG�v���Ԛ�����X����<��Q�2���c��D�·D�u�M�Ĥ�.�E'{m׎���^�?��c�B0py�Y�k.�zR��x����rS�~�����0^�WqT���K�].���K�Ql݈��
�J��Ե�-�gl92v��ܶ�
j��������\2�RD��]��\���)�or<�Ԭ�.��`@ś����2O�PF��e���n�;����"�h|�\�o7D�f�0����+s�uf\w���]a�(tAf�2%�T�l�Y�O#�l\�}�����W���30�=�E\���m:��&��0�c�D��B�nG�t��^
��Atr�q�x�6w�|2��C2�����As���t`�� +JRVb�%�z1zt�a8��z,T)23�K}���MO�-_�!�Qb/�^�Z)R�W�矰�|����Z� "��:1�ꙛ׺�����M��Ȳ�Eיj�x�<~��};C�Ev#��� �>�BS�G�?�#,�L���U����}�-���|�����h�4��2{�u�6���������`����k�s��?��H��& [ya�8�|�c�f�l�������$��E��TF6�$����#�4��8�jw-�0*Vi�?5?�j1�e�O���*F7O�5�8��o�*�]h�h�2w���zY�_Wl�1*�sׅ;�"���a�nF��1�ݟ�z4!.b?[1�$���I�y�wjV�P�2n
Os�ȉ%|G���1X��Y��<>���y���nX�,pGъ:jme�/��`/�p�D`�������F��Ā۾xߠ�QU�����<�N�w��*`}�:\���9�`�$Y��=׀y�1:O��������|�\�OG��m.�JS��0�Ѹ�u�Y���9!+\/�uO�ܝG���,k��=$u�&�0��_¯����4�'�?<�,�@Zՙ�&�ʼEN/�\\�lxtM�E��V���+|��5BHD���$��\Ȍ����V�^��v6�E��V��N��`���uE8��C�'z'Օ�&����^�3�`�ș��4^:����΅��L���m���5��Io l�/V-(�M'�a//*�D�z�D8yTfr_;�s�����Դ\eac����*`3����H9�����V�F_{����,�PE�w�u�˞���]	���hG�R!,- M�)~(�B<Jn�kk$���]4C}��Ëj��;�Y����%��6fƟ��i5�Y�΍/X���ZDe���<A��F��m:����./
%$g���z�Ab>����%Q��q]�FH�+M�f�$|� 0��,��	��\K�?���Lf���u=,:g۪�q�\�?���^�۷_��K=Q�{qW���2OF��&��4�_Py�Ŵu\S�>X�A*:���Wke�0PNޭ׶6Kv��t�(kj$�b�(w��ٯ�{�_/V6��I��ڙ��ȧqѩ�9^Z��Ti-.9��lH�?2�_Z�񐁩?�����bT<́i{��G�Į7qA�A�WR�M�}��L�S�y���Q���	�l�>��D\���# ���HK�i<^���P�
�4������ݘC�a~��.ƒ�p�w>G3D�ik���	��:�#p@8��	u���b{��w��E�e�
sI�7���O%E���"�9���Xm2}��X�ށ�bo�N��6�E�O�����;��aƮ8h�!�(켧l�9SJF����8�I⹑�+4w��jd��`x&�����Щĥry���&w���� ��"Kk=���hfQ�L���03 !�u��H�oϓ�}pj�4���M��	�������o�[jC�2$��4�w�CZ�t2�,���9~R]��Э�|!]�T�f�1=��&�e�Asw�jQ�.C�콷n�Ym[�K4��>���9 ꃅ�:��ck�)0�˳�?����/�1��ߋ�)�Ч�ǭ�����茎������q�>����KJ{1S뮤�K��j�����ji�-�1x����D���1��f�D�{�lQ��� WD�f�zS[��y�^��w�����p��F�|�^�]��Ph*�^�bs:���A�OZq��?��L|�ѥ� ]AQg�1Q$�c�#��=}�Ӈʋّ��J��@K��s�|��f�F�R;=}�:;s�Ͱ��i��$��+�r]1�~��"3,�L1�ZAe�ﰞ��%\Sb=�:��P�v@0��o��f�uZ/��/��TA} 
%ҶǊ�
�e��ԕK�@ >[J�RǭW�,r�5�77+�7�'���	Ϗ.��[������M �-�����gI;�Ϸ.���w���Sb!{}��b���� $�`ڵ�ڜ�6�W6рs�zh���Uun5����K�SZC���|�4ߍ����^l;��a?s$� >��z��	1N��y�ݓ�R7��F��[p�[cG���<7�Ƀ��Z�c�<���5�(GRۖ���A���A�9�K�*�:岞Y=�ؼ�'̜ݧ����(��Z����K��Z�uM#rV̷�w8+KzD]��P:�n�[d����;�\g��cK�}W@��x%�6@�Y!l� ��_Ug����<5ȳ�׍C�D;�Y?�6�MS��U�_�{���� 6Q�ǲ\s�p]e�v7Q��ֵ�������~�{�t��!� ��z���B}P����z�?k[|��
�y���F�z��ŧ&�̻�ZWz��X�X���lX��%��e֫��9e���������h�����搚�ž�r7�Ý:��Pr��CM,� �yV�VPt�Ie�/��|ne�h�"�����ڮ\��4�z��OJ`I��f;f�Y���,��_Jؾr@�`ꃟ�-���4
�D e+=�_�{������)Ո;"�d���ҥ{���qі��3���2Z;/[+�+ӑR�i�42\�x�����'wo�'��"˕��Isb�(���	�Rk�	[��r���/<������5��,�C�EN�
d���=r�22T|62I�A+F�!zه�yd�����T`|�l�75���a�w�&*�xKVׯC:7��cڄ�H�z������w���]D�!cR;R+6����)��ʌ�ɞ�O��uO�ZW������%oܹ�%�`��>�0q�o���3"c8�70�� �ij3��{�I�.�cZ���d-���}��خg<����V�x:b롖��`hD��bD՟�MzԎEp7eN`�,b�.$<nq.�v ���l���P*���5#�\4㩝Yn s@�^z��,5�nU'��8�1�Qz�,��;���A�*�x&H�TUTͶv��?�ʳv:��}Ɩm$,�P�X����6� ��XN������S�{�>Gs�kg�:]��Jw�9$�o�_C��\
\�!(8����S�� iUX324���2���~	zm�����m�d�� 
��/b�t\��OPs#q���R��r��O]A_����E6�h`ϗ��ˢ��a2D�&:�;\���� p��:���f�.����2�|c�g��y������je�Ͷ���3�D=@��ɇ�����3�e�#n���D��x�p-�
�L>kq���g��-n��
n��"�:ԛ7(c�c)�̋ƙ o`����lr͆�m3�b@����D�^hL���y�-j|kzA��UN�E���/Ǉ�5�_T��<��ܟ�4����sV�R�/��zB}4��:m_M��T�O����\�J`M���wg�u5�~A��U�0����s���?�R]s�d����{��p!�/�$E_�c���{�E��C-d�����N�e�$ap	�5T��Q�r��P"g�ZA�4ç�0�Qڛ<��z�臐��)��k���]�����f���T�z�92�p��ub����
�/�+��G���׹�b.~������o閅!���<kN�>0]�sKU:u&_���sF��|)��T��L�sV�Kj@�J�_`!��Σ�����G�,�>F�
.�~I��|v�â~���O�ʜ�?������1��7�TV�*+�� �)hj��Y����?�>)a�E: ��ܛ�'�h~u��ˀ�)�o��T���AՇ�/�5{��p3� u���L)'�z��$�4�4���R]���Hۆ�X>})F�R��]oR��/�d��T�׏�zs��k~�'����L}]��Jq,�3�N$d|�л��a�������@�8p��
�������j�P����Y/Ә��9��V��EP�����r� �R��R�@��[CTD��N^E.��!���㕡�����pJ;��;[:ў~i;S
%���/i�4���t���(�yI�/b��r����E@�,�CbTK�IT{��Ɔ�'{pz��:���p���g�h�^�٩�y�*�������!���X�K�Wؐ�^W����K��!�����:ӟb�&�$����� ���a�⻌(�n���{F�s+�elW2��]��4��u�����Ұ��<�P�����  �Z٣Hs-������A���]�x�����J�Y���n��`���iQ[}�]*��z�7��2�Qp�ķ��=�q�t�Ht��9�/��v������(e�X
JA��P��fj�u�\j��/���g���H+AuT3dk/�L�t�4'u���������"��л��'g_}����M8)�pe�F5�����#ֱ:V;3�KGK?ٶO�g���9cs9���	�膎�3\ՕȮn�Թٍ��˶?�ȴ��g̲$�SA����-^`���j��U���@�����KԢ�g�p�q�w��h��ɿJx�_ہ�to�j�%�!H֐5���E����{�.�٥�f��^��T|� (�)��U����"FA�8i$��:�d�{%���f�P�("��2/����$����p�8�^��4m�v9R���檪��j�[_�~��Г�~ؾl�'�Z>f.463GӁy1)��o���p�ch�����?#�ō�#?G�w�=B�h��~S�UH.µ�T�Nj���u��^J*{crN��
#���=��&j�����	�T-��^	�~"S.|��?�S"�5)l5hsȻ��n�LV�"B�9�^���w��0�p@X�L����L�������S�x��w�ºY2v�<G��i�^ñ�H��(K��~G�d���a��W򽲺���Xֲ�ؤ�.P1տ'���Vuf�y�+��s>y(}ơɀ�I/O���e������承��Ѕz�}�U�`ܹ��{�����/�|ַ'�j�"���K�� �BI��
C�j�*>pf�P�9d����@�oOR��=��v%�s";@ٔua�4�_T�G�%d����iٳ��;;�$SK�2kwi���o6���^��s���_PT)��la��Dȥsd����}R�-++%�+ޘK�7�I�VnQϞ���>bP}&�5;�	9v�h�wO�d�$~��xg$� ��������I��*^=�Mw�v�T�ex�?�d�4rL�iǂ��I��?
�2G��#|�d���S$�ki�r�!�Bs��2�1J[#�O�/�'8hbx�|K%O�23K�����_U������(+^����Z�U��S�Hn�-Gl6�^<>�1��W5�}p�ރ��K������"�WhA������9C���0��/v�h��X
po�U�p-��j7a6��z�=����?!Xy��ivyV3c��P����H�L��.�)���[�Y������L�W:���h1��-t�e���O؏9k��lp�6I�g[�_R\�G5�ն&����Ż�9�Ӆ����t�ٶ� �V������7>b��%=Dܑ)g���븬�iޢqʓ��kӜ}��J�r��H��$���[��-+Ks�ތV#�o�����|#]���?q{��������E�r�,-�M�vv� r`_2���ƩQ+I$n\����4��{1=K�Ԃ���D��\�7�����(m��ܝ>X�7u�����^��.|�,���#x�v-�)���&x���8;�t�B�ɮ?�=s���:�`�qV����T�\}���V����VvG��BMO����}h�R'�-+}9n@�R�lY8��]	Vh�3#f�0����aż���vY�JJ@�C�
u�Q�p����֭��
��wS�[1�������b ޢđQ&ë��v͒zhjH�N�t^ִ�Қ�x�;"2�E�jP+Dg�4"lܪ�';pZԉ9/פ4���;�HE/� "8�oݭjf��1�cP0�l����-�3|5Wit��Aܟ1��\���y���P�Ѕ2����1�r{"X��Ľ��D�=ZҶ����&UD�nQ���;C�6"V��UY��ۓ�L���4y���_<����~�H��U��;s��6�@�*s[����l�����"�? ��rO]x�	�{�����.�s�E|�,x�f�M�K��Hzӹ�w��7����V�x@ic�f���$�4�2��-�=ۭp�6���@׹��V�g��?�-p?����q��ƚXMkrE��_kC����p␫�4:�˛W�P�݇�8��0(�w�P �����=���-rd�����=.����dpfr���toř@҅�(�l�~���-�X`��9�ࣾ�Q���G��3�}��-�S��W��EHu��u< ��6�-���m�Q��}��z�4p9XyP`�&S�w�b�2�e��^YQ��T5�����Ҿ�C�X(4D;�o���/��Wq{������:�x�?��d���t�ے+�L�9���=P��*�X�hmH�Zq��M���{�A��e�א�����\���R�p�<�48�M%O�aN��ļ$H\��&��ɟ�L��h�F:,F�a44��?Q�Wb�}/8��+�P�G_B���e�F������L�N�	����fc���������ל
N�g�/<�t����:he����Kǹh������bf�Y80�4��<Yu,.zJ�qy�q��H��~f���8v�ѓ~|I��#�6������<��+u�/�����)�=[G���,`0]�Є�U��XنS� U��3`�v6X��]��?�fk���L
<��z��t��E-+�7^��~�i�r�~��W~�3^U;Y�;��[0�s��8"�3c��Y��8�|T7����X.�E+4O����r���SK��Y�����_�й,=h��@�Ы�9�n�uP�21>�*�65+�6ׄW��e��K��Vx����� �W�+�m:�����[,c�g%4q{�l:�P��
ټ1�<����2�R��璫N|o"j�/H�7��x1�U��$ȉ4` �B�;^9uo�@6@�����__Q�m��"ʬh_�7��|	c-L��l���v}�*����i��j��^�0G~�\Dkm�O�\_m�q����jjR5�L!��5(C�{�Af�~��}FGerҒ�+�)t^�\�`E�XCһ Q����y�,ԣ/v����h�yǴ�Z�׹;�p���2�sv�^�������trԠ-�����<;��|�-�S�3g�#�E���y[İYć���۽_��r�9TSo��O�ׂ&zQZ��"�"ժ4�6�	�;�ރ�f!ìe+'�/��Y�#�[3�w��������qG��Lu�5�4$�!���,��~4��{�L�Ҋ�`
� kO5������aE 7���w��G���م�}]J�?k�Aƥ��\ԬN��3��!��JB�6�I��,a��!rDݍ
������Vm��(I*Ì�c����j�V�η��%�ΣC�0B��������o��.�n�*c�F����g2>MU��1��9z)�ڷ^��yT���"�vG]tS�Խ�|�#��'��{�"�~{K�S���l�����J�� L1ш
�T%���W�j��9�#��������%&��)(�f���{��ƅ��(
b~�@3�f�)d4����Tl�w9X�ຏb��H����ԓi|r�UgtGq�҂�ow�)���+�2i��[�����AMbʐ#�8V@��Aq�36��}H����Gx�,m¶jא�2����A�]���uv�0�Ո%����:5�F9�oų�����9�JG�R�+ۙr��/��e�� Xp���\��J���k��	��Q�a`<��䢹*�a���mM y܀���jGC���}�X� i�
��E��? b,V6��Tc`�X#:���O;��_�c��j�e����:!IuK�c�'�M,��\��,,0qǺ?� e$_��Tt¢�{;*����LG��~w�&�!oR��z�W�*r�+Tk���]�s.���OJ���!�_�΍TX�E
������j����+?���Q���P����/3-3mhY#�*�Pb�ڪGy)�����`|��y�\|3��V��Ɋ�ߨm��x�sz�P)���I/���<�3�W؟;RZ3Kz�}��J�@�`�R��_��V�I��P]6���a.4y?�� �G괍�;9xu/��g?M�����k�XWB���}�Mh��c���[a�ͥK��n�˗ҫU�����6���O~���{�,E�tٺ��z���V��M��I�P[�ֽ��1]������i��y-�p>���qYp���o+9ڻ]*i�oe�M<�����������Z%�Ə�R%[;Y��d~(S�ʊ��L$86�cߊ�	]�D�D�����r��/�u~q KE����!#��6p�u��C�xM,����X��~ְ�T����e9�3>-��Yi��ȷ}�1�m�f�pNu^�ߌ��6@��c��E�>��?D �ͳ~�a�Ѭ{��qN�ښ��yЍ�8��^=ew��m�����r}�^8�~��ʷ���g���U�vyl���z�×+,1ձ4.�k�y����n�4e4�hcWd|�Q]ͅ����2�S.��%�xy�rk�p!/�hk�H�ե:v���ݫ��/�����r]��yn1��ͺ;k���/A��.�n����H��>u�	����da�T�Tf.��A�D�l"7�0 nW�}w�ا"g3�W�h�5�YXC��;f@=bC��.�����%ғ#���p辨�Cgs�Jy�;ccZk>�ݹ���������0��Ϥ�� 9�r�:~=~���ș�۲�P�<�G��F.K�%l����;6*��X�n�<��ӼDq2�q�%��ma]���/N1�˸�����tFh��- 4���v	���n�h�ڡj�*@ J�iO�������y�uwFΣ�!=V�"�i����V�c�:9tT��3�fu Ze�s��o8����1rf@1����	���]�!������M2֚d�%O����ؽp%�������I���+���j>��A2~aǥ;k�d����s[]H�eB��S��2T��#��O���2��ʠ�%R���՛���06��e���ڼ	��gW�"4�A�)�L�>���GнD�_F�����m�~܄����\>ggE5R�b�g�׶|��,�Q��ó��[�6���'K2���;���dP�}���n���&�=����Ͽx*<��f�j���C���DW�kV&��&�������V#�Ŝ�Ƨ�ߓ�j�������?4�D�
%���i�:�H��ͱwI��̌��}��(��<86�qp�=��z�������yy�s����������Ih����؜�5Ts7��+�ag�5tg?�DN����z�:;��;�\��p���pg�G5NAA�[5�/c�Z�_10<�u������Y��7O�~�d�����1��e���A���kK�[�]�c����g.���B34�xa�3��j���!2b�����t޽EG��}w�L�z�׻]�#-�r)�����.k����r�ůN,�������;���>�-I^} S��5��x��9��ڴW:@sv
Ch�w}�b�D ����x�Ǎ��a��\�n^���	�Q)\r�cx���2DAǾ^����g{Gw8*�����Wsv,'�r:[��zw�����Р����t��� a��ƞ����?�[��V�Ӹ��S.$Qs�1�벍�U�UA"G_0��8��+Y���������xB���/Ϟ��+�ˍ��:��>w������Ċ�D��ٝ����˥|����6�K5|=��v��Y&e�����?o�J��͟��s��\�q�ፗ���X�R���n0V	��srr��~����/��( ��ttha�M)s���.�ݻ�)��s&%��)!$L���|�䮴�j�Z��3"n<R����$������E��`�f��t�����o�x쎛o��Z�'��>㶱�'��C�b`�������6/d�F�1�53m&A��y�L��k>S3�\�g��յqV��I�9}`&��_]�. CDz��e%�w~r(e��L����?��� Z����s�o�Pf���)&
����.�4E��������H{��v$��I�M��;�1{}3�����De��k5��F9�\h�e�r��H$�d�\V�C��صۤ�<��|g��Ե��ū��,���
�=)�����=L"��b~`�r���Eh;=!�������8'5sʕa�0�1.�%�_����d�H_ji�~�`qRs��ʚ�8���}	q�+uU|��W�����Ş��E��e-�E1�]-���#J���R�'�6o�/�����ŝ6^��K���$�_V7��P�ѣƈ�uО3���ԑlu��I|^��N��7X[���HR��!��t�2m�^�������F~��]Ж���g��~Z�M����5�����~" 5'V/w��ݟ1��\l;	I8� Ia������a�I��k]6ET?�lm>0�ҡ[%�|Ԉ��.�q�^[N��R��F5��U����H"E��<���Փt��O�]�f0���{�%���>���/{�u�0�Kq&(HƢ`�o#�!FX�L���tV���F�Z`��H������9~�hSb9o}Tv���8DA��진����:a���>*���>�E8R�����w �5}��l�U�P;+�1d�;-�wњ<#�'�t׺;vI16��4�F�y��.`���Ţ�����Y��h�7B���7��(Q�d�u}e��e��R�1�ˑ��Sn�f^���u�~}����^���le�Ϻ+�VR����ɣ��%�s�]i)�Ӧ�J0���d���or`� ��ӌ6�#��޶�pk�����cآzx?��K����*uG�{�^0L�F5=^#~�g����%�%���RO{�=�����6�g^�z���țg:zӮ4�|�'>�\���|#�@~��G���y����z���t�� ����+��U�ʾ����,�}_^hI��fAw*���d���L����^>Y������=�J����;{BJC�S��M������Vo��ˬ�k�"�#�$?6�c߈l.%Es�ю-�	�<����3Ō�i��OX�� �b̦�k�6m��΄�+كA��������yp�/�R�Č\�.u�+�������W�ޙ��7:/��3�������J��)�/�-���PP Z'W,ǫ)6Z�?!
�y��I����7XX71���1���_�,�j�ۺf�"뷓$	��=	6�s/�ow�^��Խ{%kV�93%�#�dA�QN���$.n{$��+��Y�X�BD����bؖ?6�X{'׌ٝ�@�8���Ɏ��GU% ��r���*���2Tִ��-���5��n����=��K��dϝp��[N-�	f,�YG�d����f\GyY�|��}Z����[�	�A��E~�a��m�O}����3�*����d]՜� ��;V��nɸ�IFe��C��݂\&� @�E5�}VE6{!M�'�����/v�40ޣy��[���E+�_�~P��E����L�}��1ڲ������Zڸ}ݍ��n���3 DZ�9^ƽ=k���VK��]��J�,f1Kđ�;��;��h�&��'��q��d ����9v�%���
�pj����?4G�~��#���������K�&H9P��y�,y�*��Kd��}�U)�z��7�2k%!Df���Wc�{�Y|���ͫ��G��F�b�]�����Ri�4g��]^�I	�j@��-3J���)FΙ�Y2�E�1�K;�M����:�Y�W涘�ؑmCO\;���zeu��X��?pLs�~�H��{�-{^T �s��z����j%# �&�;�����!��l78����L\b�B��B�M�g�_��J,[~Y=���̢U�S6p)K����K��_Ӷ�eX��O�ןii���-���7������&2}��K���Y.���p�$9�/��Ϯ%��E��qfC^��K���T�@�I|������_ ��y�C�rk��`X������Zե��L�k��y��HW���Bv��������fh^�ĥ�BRg�	�#ll�F;����w��֍i�F�7����^�
���jq�[��7��륙v*Q́<��ka�/ɐ�'r��=�p�l=k����*� /r��ŶÞ�,2�� ���e���U@��^�k����)̣ ���{G�|Um��]�
��
=�m��R�i8�����H���Y~��c
�H��.e�5o�$���f���*��0l��(�Y�_IH��,�i!�A��Ė�(ՀΣ�PV{>�uGe.t�.�p�e�� ��;J���$#lY������3 l����">˂�z�ێ��曟G&x�#I�N����I���G�N����#��D}3q�B���X��{/�G��VGb���ϛ�Q�u݂���w<;Av��
 ��z�V<3�� 8&j���^xV�Sf\�ڐ�����zJ6����;��+���� ��X�!^} J�;�4xy	[��Ks)�k��<��� #-`ׯ���3`�cvD��/ܗ�]~��*��X�8ſ�*aT�=6 �
�:gn�cDc*2�T������l�]Z�"�$�e����i���e����nBTnod�߀����: @����\�s���?�4�D�Lu�*�ML���v82�?��R�C;���O����Bj���hۿ��HK['�2�σBv;�m����W�A?P⒒��r>�a�k�?��9p
�6�UK���h�t�����TzM&�{a�/\_0�����%�����H�x��P�&��OM���Yne1�X��9��Ul2vCC|I.�r�n��^�7��4N6�Q
�Xo	`����m��@\Q�5�5[�U��j?�zc�"�[���V�A�Ǣ,Ⱥ^}��������L���1�.�o1[�K)~��°I���e>�9�F��Y�3���)= +u}�b�fW�cw?l�6_ ����/ӿ� �
"�]�?�R�v������	^�
��	�9�^4.�B�l���X�~;��\�N���x%������B�Q�b�m	�#�9�X��[D��֞��S�C]�6�[����}F��7�
^�~o�m��6���/�`�ce�%�oȳ*։����~�����Qp?JL�Ϗ�V�x'-r �W�xU�?^�~��D8Qp&`)'O��1}��ȷ6*r�J�����yB�P���ݎ��g*�d�4��\�����Ù���B���]F_}P��N�/.����6��
��K�f��j�
ܵ$��tzͲ����@J�fvX��Y��hYT�t_��Qu�� k�L���ӣ��	g<�JIBա���O�II�{tb�؞̜��[���4�Bo¿Z�'{*2&�A�ǐB5��P�z��ͭV�H^RakN*�I�F�<Z�CY�M��t��W�~�Onk~�|�~.���|n��Ni�6��5d�cu��v��|���VL;1	Q{��fz"H����\F�Q�P6�����Q��/��������u�?�9�L$\{�Aʢ�<$�\�=M��tk�Spd�0G���	�.����[�LՒ��8������Q˙;��?y�0�m�|��4��B�3��qgG���'����Ŷ�,�$Z̽)FYVf�/��dg�D�q8@�kn���KRB�T=�Ӟ�}���Qn|N���~��2F1b�)@�o���+��{2o�H��4Oka�)��ҷ�:!��ڄկL�b�@�8%�� ��}��+>��m�$Һ��S�H��p�Xw#�
h� ���o<���u,�`7�Ze�m���q�{��;]m>H���A4���~�0����BMy1���U95��knU�R�]L�O��������V�)��)����������̠b�"�_���-�_
U��I��P��EP��ʹ�er 	1��C��sv�����-Uk��Mk���d��ۙW�oק�[祀��Qd=���GbR@8�uZ�P�4���+�qV��Vv���lP�A&O���9}F�%j����'A|Q+�.�	�;Z�rDBc���F��SI[��I�r�^mL��^8���sw4��7�����(a���"יF��\��b�+W;�w�"���e-wF��3��0D��f�g9W�a]�y����9\uv�O����Z�Ք ����{�t+�A>�T ��J�46'��.X�[���12���g��DW�,q�Y�OI�qVh���:�������㎔ ����d_�;�'�v7�m�4����y�����M>�x|����~��������
��F`cr'M(�*+��ŷQ��!�K n���N�D�Ԣ.�'��������JA��T�G�$Aܞj(�� "�*����n�>�����l��-r`�����HGl���OƯw�6��{yG���ҋ����^B�����g����ۡ�3��h�7�R$8y�K�*K�il�����A�д�,����`�jM)@�|�K��z
��В���B�Q�������sk����n޽�k�3�
��Dep����cb��}]o��^����Y�x~5�a�ViIH�Z�\��^2��3{�t�>�fU[��^˱�b����{��a_��U�b����ʘ-�)�84��a4�����Sde��Lqw��S{=d?s=�ͳ���U��S��P]��k%�Au­�:\�ˬ;6R�l���I����.P�ة�L������cI����FF��'Ԗ������*�vܢ;P��3j�M��B��F ��I�mOq?���0�A߹WП3j�#QF�n���(ն�l�q�E���s]��!��<��6�I��$eU�l����D	�'�{win6�ao�H]o�X��]H���"#uN3���X`?6��
��9:�ڹ����1��(B��~��M�d�^�R��������%��B�d��2����3��@��Ȃ>�V݃JJ��v���8fV~���Gv"��'��O<�_8�P�ҫ9��;�u^H>�N��I+��ꂎ滬��3˱���V~	��p�h:%�|�����N?�2�5����鍊Ur.�]	͐>�I��3��j�y��s���{�3�/�V�����z���Em��m��H��o��B�)��s���KY��d>��"�d��u�����cS�(�0K�*|k�\����t*]�Kg�x�����7����7�4�v1�4Q	B�����H��|>x؂�)~���	.7�?��,�{��e��ކ7��]�u�PF�b����G۪uK9�S����)Q���ن\]g��O�2�;h ����ǘ���7�����v� ދ�])ǋ%v�
�]"Z�ΰx��f� ��� �g�Պ:-��rYa�E�,��>������'���j�I�~��Em�w��)��Ÿk
EC^���������F /Ȁ:&���h�r�CinŐ?� �����)��j
����SO�+�-�����'	=�� s����q����r�U�)�n	;��ƠH�
�a|2 Pa����-���AϬZ�N&܈[[��?�bTb�i*x�~\ga� T��Y/|�zc$��C��g����������������2tK�3l�W� W0�]pS�K(��T�!I�)�������Qs�l��<G����5b�d�`��yB;)�NM: �7}������^�6Syq.FGJB魌�%�?,����F�vT�F��0���=�a3���<Xqb��DR�� ����pl�q�ٱR�~�m�T[2-�l�)��D7[6���B�Op��v�"Vs.�6��ڽ�N<������^��K2�⋢�GJ{��e���@�pZג�
�-ʗ#�8����d��r���@q�]�}BgOq���!�r -�pu<��< ��z���#�N�.�ur�p���Z[�~a3�;3r�X��L��:W�U#��I[��ל�uW��7����{��;'���zN�闕�6s3~��WG��v���p��Wb��`�V籾ѣ�p�L��xx��` 6��A`L�/r��X�*���RJ�b��������)?=p�6�������gM�G�\MσS3����#l|[k�~���.z8 �?��-Q�'m��_	4>�/�s�Z� � ��u6n~ݱ�z����i�iq�0��{�t�lb(�ނ�E�&��;��Z�XkɌxuEV�h	e&<M,�CMm9[F	8�r�Ri��H�Vk�Xa� �YPj-(!+M_��S7�u%�@5�`��Yz�̕��=3�si26������g����d����u�b	��Reyu��7�+ZXV�Tu�фs�m!�f��0O]��7�L���������Cq��_��>���4�8*�3v�-ɮFE1+�/R���[ꐆ2�i�m�m(�
��ߑÞa���yc��&��o�K&C��-*:&1%��@�,���ʥCsݻ��q=
x:�نo��/�\�!�?�ĭ��H+N�KӃ�Rz� ����E�!��l����s�v�q��Z5�.ٴ�?s����F$��N�7�-�HM�p�T�*�^�����xp���.�/O9G[ڴ�XP���IIT��s���X����䱒u�f\	��o��أ�W'�2�S��H��v��f]�t�,7R��	x���E0�9��_��[������PK��;Q[F����n�<-g`���!,����U�w�����E���E3D�NmS�{S��[�P;%u$:::3Љ@��VV��J5���+=�]v���։�J~	��a���{�ݳ��g�d�b��P��dO�X�~�p�SP���#�&��LF�_���=ܣʑ?�Ԕ|�[�'�})%�_�V�KY����D�����{C5nm�+��X���	R��@���ݮ	~d�U^�s�?�>{K�v!��0����%����	��k�mlŤ������n{�g9?�$||��r�����/A��(�s\!��K����#c�v�P��Z��(o-{��V�5��*1�������!o�(�I�T������W�8�&=_c&P��)<u�J�ݍ����� �05	������$a��Uq��� y�Ι�c�g�M�
:=7;��6CgJ	�C ��U{�U����%]��W�D)`��>�|^�F��(�k� |m�(����:�<5mpa^m��ă�1�n��ۊ�R��bS�}0'W��fZ��{������:�����O��2�	���-i���=|&RL|�����k0r'桲^���{�b����|ANe�際��|��A��<q� ��.���1
x�t�-�v}6���6wУ}���=3{���%S�ly��  |��҃U�%�bߢ��%�7'*����umlA��~t�� ��	�-�R*w��ݤ��g�}�iv��u���7ze�������y<���ڀ���֚ٲ�&�^>��I4�чN-� ޑ����YI��ұ�5�hAe���T�����P5�>�e���j���3+�>Z��4��>���oQNO�$�bG���%�/j���ÿ��	Ö�QN��X?8������*�}tj]Tv�"��;L�Uf����/?\>u����C���%-f3����^���ove��`7���o����3z����E����h���E��}�&))��m�lREm�}Է�3wx�X2�Pf��7=Ϸk?d]�H�	���;#���Sb=�ռ���?�A@��Yd��^��JM�8��Ҁ�^TD|�s����1�� ߏ���M�۝؟���K���ހ��v��}��/.���Ư썯��b�qVU�����3�T����7�h"�깂Ȓm�V���WdHZ�0��;C���u���x�%64�o�'���m��Ύ�x$Y�����q؅q }���8-�F��$6����'�<�j�l��}"OK�EM���;��ڢe�����ռJR���5��9�&q{ռ��=�E�c�!�  ���Z�ZQw���A�n�7	X@	����9PK/�;��QȻm�0��K)\3����W���A|2�	�";��p��_g�	THS����_o� ⍢k�.t�eV}M�����n��}|��^X�OM%n���KdM2c���>��t�ީT�]L�g���r��5�|��zk��D�p��<��(f�N4Qi,b'Z���J����,����(;�Mhq��ȑ�$h+�0�G�'��k���["5�l:��`{R��ۯ��X��y�7�����S�P�c�I͉��-4�b���ƹ�ȉs2"�o�څ�y����
 ��[UBM~���wO�@{)͆άG���Tx�����xN
��������_���I�C��]�
�~=d��A�[m]����]Qh�������w��,�'����t�@�t���H�j#{�ٯ�k��[�ڒ �2�h"�e�a��PG�qD�l��(�����zN)c?�:��|�T;��H3;�R,T�(g3�w[{��?^\hU��ɒ�]���ݾ��Q �z���b7��F����|5���{� l���q������~�L]��<���.	�t�/L���gj��۹�jTt6��^f��,�_�x�M�_��wXO��vx��= ����;���w��P����aP���+��:0JۑC�}t�a��h�h���Wmվ��s��{�-�{�n/����c��6Va+��E>���3$-�C��>U��p��ܠ��0#!�c��o�4iq�2MBlO#a7j��D��ɋ��!
?P���U��ޓ'JX��%��NA�B�<���#u6ǧU-mSܪu�K��ǂ|�
6�?kt�������*鬒�}W�o��uxz�����2)g�5fi�*	 ?���fK5��E��Y=��k�Tg|�*̬�</��I@!�lzch��zE�)�M�v_T�4X�
�"C�}�D6��q�dBʹ��7D�{W~	B� q���G�E~�>/ľUk��}yƊ�xBQ
B�a���n}����s����}�l\P@�䟻\q@�خ9�ފ@!=�l��=�F2����Q/2�;����p����4]}�d��To��ο��r���yɧ)��7��,w�n���?�/n �.�k0��,@��i��kkqF��t�@\.v+AE~�
�F�:R�9,��0��~"�	8{��+��!�����_$�{�`]"�#�
��Pio�]��a�+��Gߑ�󍲍�E�>>��	xjo�Z��|�@@XU�P��Iׄ,0�����߽��d,�d��Z%(I���E���$�!�� �p��@�Ŷg=����Vi���H��mv�>�N�lE���_��X��?4(�����_���$��2����S��gǽ�4�:�d�X�ъ�7B�g��r8�(�	�}�GF(�e=�F�h���_�/�s���)m��"~Sz�|�$�<�?%2@<�����e�b,=��ae:��d�q���zY<7�����=|��WK�X��{��~�jSa�L6a/����a�N�Ժi���d\��^�'�����iJ���80�����}[�H�a3p���3fȮ���8c�8�7�},���'"u��V�d9�Z�o��^^{u.��^�ӖP��Q%��������6λSR�Kr�/��E��Q|��ْ:���g_/��^����?���3�5b�K"q��$���lU�7���w	`��k�wcǤ14���]���3�+1 r�t�xQƿ�q~Z�[P���?�K�ah��6`զ-���}�O�Ό����4"��UW:�!f�Z���z�j�&�wQu�r�Q	�ƣ���&.�%��,8��Й�_�&�e�|�ִk1=lμ@�x&/�_Os������8�T�BČ:��cn�{��\d�:M�	ʕ�uj��̅ v~&_N��g�����)"��QP�x<x!k9���<Q^�w��$22B�+Yeyj�E��n�~*�D�
��S�M�1�4ҷ�I3����U��Xɾ�c-^Z����������2���8���T�V��Im\.��S�m��!��}��!yO�(v-����z|��*F����T�{W�����H�_��
7�}�Z"�v��+�ry>�H����Ǚ��/Z؜vD.Kw�~��}kP"��� ����b���t��R���0��B�$�܌X�J�&\����]Ș��@�X��z���}��:1O�$a ��Û�����7K�-��[a+������nnIj�~����N;��xȱ�~�{p?�:w�a�����5�`_	ܙ~ܱ�}�J�����ј��df�4ѹ5d�mÌ��7t�0�;�謹�%�2l�YN;��|��J��N�T�u���!������s���/��������mw���iݗ�����b�a?!x�w��p:�r^j�3ߑ�'8�1:�e@���y��������a�s�_K���*̟����x]Y�F��#}�a�݇���]��צ�Ȯ#Yڝ�m\��&r�-ܿ8�e�m	��Y*�$��Y��-W*{�d�y	��_��2`��su���>�/}F�� 6�V5 G��ݛ �8�3�Bs�#v��	j ~Z�1xC&�?�������-K����V&��+''O�!4���b⪪�R�*?5��#FFF�R'�)����]V���[��\t�
����χ�v��	RT�Aܓ��ư�H}�L�:?X@��_�_���t ܊�����~�/S8�l�Fz-�{ߞW�P��3�F�ib����p�v��Þ��6��A�WE�<Ӽ�=��C��!�ã�Ͻ���|�����|�ɜ,�{5O�%T�j��5M�z4V,$��/,�.D��3�.$G�Z,ʣ�sg���)����n��H�p�%��������hF��p_���n�Ec�R�AJ`�HF3�`�Vt_]=2x̧�+�e�U�JZ�>�o����W`<��]� ��Eʿȓ�0�QvTECu~C-Qb�DE���v�@���9�<-��2��/���Xө?PJN6S_>�F���+}����TsՂJ��]�ꖏ�Ph��CJi�����v���Wd���"+�	-�GX
���ƦyQ�v�;9�]v�	��nr���b�Ž�C����Vt��W�$�gk�UR�Ap�>�;�K�[���{?���?Ò�n+���vQ93�����:�J���s�姶Ս���4��>��'����~�jȽ�	��Ʒ�9ʚ�����F��������g8�_��~GQ%�Nm!I l	N�B�D�Y����/h|l���e����۱�X��8�`��W��8z��]��PO�xo��A^�o;F���]��8o��{�M��r" ��
�^��j(i7ij�x��.ד,����Uj(�Ĺ��������3�P�y�_CV�5=|�YqKP���+�B�4����-�J��V~�] u�ȖAd�,q�C<��#`SWBD9~�`L?8Ǫ�V��%��'=LW�|�M@�M�꾴v�M�l�͛A2���|��][����(�f
�hLЀ�5���{6"�����1��F��t#��+n
�f���̓E���{[�`0�W9�ʌ] =��4�%�<���d�L����ƃ��2�ܹ6��<� R�e��x�B��[�4�a�E����o��j����:�h��%��枤$<��)��=�=���)�~;��O5*U	r��kwP4�$?��"m�'i]��.��������B�4_�hau�Ab6�a ���3(1Ќ�X&�Z�����w;a<z����H\� �6,Sk�m��φ竷��`�Ó��#���V�*�����yt����V��e��'�0P�\	�������F��u]m*��2R��
}ΐ{�z���t��UuB�Y/���!��5I4k	����
�-�Ɩ��J���/���d�N��yA��:68l��,��ǋvWԝ�a�-��K����������|�j�}��<X��R�H3���O?��-̲���Jޣ��xW��v�hy�k�K�o=�Շ9�}����)�*�1�&l�Ÿ�����"�a�|�X<&��%�G9���s�+ 6�-�E@��gaoZ��j0��/�����5��E�����)9�Hɖ�e��\j��V�9�� E���ۑ�ܽ�6n<�ê߂�70�V��ȶ�A�Wr�V.���%f����]�U��tV���/{�+�Sa\�7�VE����� �$��y��c����A�xL�v��q�yD��J�h@Ր�&]A�`�HeR�(��#��<��R��Yϗ��>����"H�Yֺ�/`�0/�QZ!!5-����jBO>��%w�ZD��K�(��r��dJ�}d'ڣ�f�pg�~E�o�o	H-�|ض�����=S�̦��B[,���u����k��g�>�G8��.t@�l���� �C|��i.=&�����������IW*����!O�U.���E^�)�G��2��߷2RcITy��f�`��)tΫ:�W0+[���zxV��)����廊=H�U�C.3J
��i����)m(�04����g { rY͉���ڂ�u'@v��)��ğ¿�I>>x�k��ڮ�N/*�k�+���n�YQ���i��� ���#h`�Ek����>���N�r�J��F��������b0�<y[��
H|���(ַ�D��
Uݗt�G]� �厪�7OBઞ��,��	��z
�K.�\B8��
��b^��|M�Hj=n���>FC��l�!D�!��#��0"��?��O1Qa^����|V솫����#�ă]��>�������J�"'�e�{` �#̇���"�S83S|�d7%�����kwP�L�1�Uyd姖�/�9���\�1�<;�H�ϋ2z�]��gx(=����Ί>A��!�9-.9�>�$khht�"�vd�-�W9�W�E�</�g���m5�w��c���SS(=�agof0�=�|��G�4l��z>��%: {�1ꖝe�G��T�P|��	~�/��
հ'F�h耈v� ����k���4��W[c�g�(eΎ��o��On>T�8�"�W��k6���V�/50-':�t��U��>�O�����M�y���?̟+�l��oO7�J��0�2:����SN_e����fx��	�kN�P K�w�0j\�-���2�O�Y��#�X�d����}�^��ЯIC;sʶ���E������)�� Ff\O�g|���,Ԯ��f��=����zqT>��W�����-�5/�ڴ/>-��cg�%dx��4+��J��e+���[^a!��4׭�����(���s�{�����Ty䥖
ڱ�h���"����2RLm˗�4�[�~M:��;˧JZ_�`�a�H͔e�:��>��F21�[ah:U�Hj�Čn���*����ۚ7w�Ha�6�YqY6K|(��CL��r1���r�9�$�`k8����i�ûMx�<��o�@L;sl�	�T�_v������=<'4��j�)Ty�����Ɋ�-��ydg:	�^����-?:�h�z���0ju =f���jf��7v����0~��5��t��XZl��t	kQ����F���w�ʷ�9����헢���^x��s�|
v�b�O�N@�N�Z�<�������f���?H�]!���ZZA���9v�����,�Gs��ƞ+��t��Q�>|�v��}�u�y�R�PJ_'1�l9Le����BWx)Br�~-v��6���im-9,@�������Ūs�ڼr���/O��>�{�{��x[��hxL�aw���_���ƽ��, ��㕄$��L���T�3\�YO���/9��ڗc�*%���������;)ԡ�!��K���q) ��Ln$�50ā�?���u(bԋFٰ8q�r(��B�����#4�Ǝ�U��Oz!��Q��'e���慣��a�������5��.�
T?�v|�t��S+(��Ī1H��T3���s<�ۏ���|QkU� �N�a+��c�M���^0��w��n�y?���N��m},ڲ+1�/�u�@��H��
)Ap݁#ӑ��l�<��ph��U��{
����R z�x���]{�'=���&�8�X\tW�V\;�X2x1����]d�d9���I%U�9��a�[�M����[�.B��_9����h7�
�����+����J�{�A�͆q\��(��k�_�U\c�$�/0@��ͬ�c�:q����7��ܢr�����4�z�a�P���?�]�ɳ����,�3�	�|=-4���q����V�� ֭��*����7p���74by�_�+����{r�}|+�:���H�������=�aU¡�[s]������ʂ�{y?�F�B��]�w��5P3R?ɷI5O�/%���jnuV� q�u��ݝ�b�.a�M�"9��_����֧>v]�#�?�X{A�|�E�����7��RJ"E��WC�-_�*B��F��K��������N04P�	y��d����}�u�ڿ��^Um�x�U�2Z���4�}��\�t�	���JT��>O� ��ܔ(�f�y�>b�U@Im.�!�+����b�����Ч������n(}L�z��]i�D��}��A���2��5�>�PQc"���
����/Qt1���	,�t4O:�6OG6?u��噸5c�'���3=�k(�P����i�~����K�i��$�k�Q��&_H(��>�1�/����w/ m�,�$���k�Pm�|�����T�;БJ��=�G�*C7���	Z[?��|[�g2���+����3Li���P��p��_���4-��|�Wq�r�� ��G��IQ��5�^n�є��5��Sd`��)���\��h��^r�$�0���q1�z(O��L}·�$7���6�0G��r�_o��3Q�=Z�󢈎v#�"���4M��A%���z��aJ�*-�u���ˉn0Rۗ�v��#�j���_6N9V2��H�8�ܟhK�.�G��Xq���?}�K�,�h��0?���4/R��c��p6��)m󏘔ЏkM��5KD������gE�EKþ4��y��ۮ��=b:7v���2�[��'֒Z" ���c���E[G��9n�=�;�}��nb��d��]�f�A�f�f���^�O��:�~6����a����P���	D��_L��_�H<�i;(
{o�U���{�vm�4׋]�?��veg�����	kkY�GWﲖݚ!�{�n=��YO�W���Se�׳�?����A��S�#�R+E���WA���C�5)��+��q�����[��>�us����ɚ�0�K[iqZV�i�"��E_饯�V���e��-+}�N蘯���mz�Ū�ܜ�s� ������D�}S�K�?5c~Ʋ#y~�G-W�q��Hv�j�&c2j�����`2�h51��I�#��&?��;Y�yH.f[��g�8�h���1���w=��'�n��Fpz���� f��[��G{�o�����]ܫ���7�_#�n��_������m�iTӥ��6ґ��]V���%���n�#/,I�CQ���t6��XN�织�0���������q��!'i����گ��PN��R��Nv��.�\�ş�q<K7�z�ͨ�\��Al��y��<:^�6욈G|u�S�4[�i����ȗ��<�������z쉙���[K���d9���9���ْ�p�J&��
��#�]�SS����g泸���&�i��_����^lEY���g���Tz� ����Q���	���ZC������L����I��N�.�m׹��<�I����)�tT���(r��W8���c��Q��Z���A[���lDS�<�& S��M*p�9�s�[�t!�:�6���5���Z����xJj;�����>� ;�l3���,Ola��:⹘QBٓ�oU����]P�}օ�j������qI<�\S]�3*)9+�΍�S��2�[Ss���A��"�1���Ʊ.�,�ԙP1��^���b�''�HsOFѬ\y ��ӵ:wZ~����.�Ӆ��Y���ad�����x��5�̟���|)�[�HaF̬d(&�'�Δ~�؝B/�C<���
��1X%&ى����s�Pjj��^�6�-������a��}���+�i����{FÜ����)gc�d�Yj�c�_驪�� b�JOI�ů�Xq�Ƽ�����~s�G�+-\��>u�>��v�(NPjO xW.5,�K�@a�5+��G�$�����>k����1�ջԚ���͋�c�{�������U�����Z�5�NꮴJ��:O�2���)�'<�iɡ���Ւ �U����a����~�.���y�`���Pg`ۯ�}�Z��v����5�B1%��Z�ym�q���s3ݓ1�I6/�����FI^��,u#�v㫋|Qn���;$�Ǣ;Tsa�e×��e��C�y����O�hL��h���Q�	�V�U��>ٛ:�9sug*;� ��T�bD�O	��e�-}���
ȅk�����Sj+���5�D~0�?UIU�����mo�y(�s��*	�94@�X�e������	�=$ �u�?���0Zf���6�>�YH	S�(�NJ�W���n��� ^���"8e$�`�p�j�|�n�d���+�_�v�f٣�G���A�C�ȗ>�s����:'*��1���t��T�ߟT>��T��WȼVY!TY��5��+Y!$d\{˾���Y�ko�����|���T��=��9�y���:��MK�����5�ڹ,�rGj�[VS�+ђCX`t��i�V�JZi��d�
�G��g��B<�{d�G�
R��UmU�D�v�]���??ml�5�X8�9�J���KU�No�=���1��K�ڴ���l�W�d
ͬ��Qe�P0��4��\h��h���B6�Y"��'�8�����r�V	�uG�������E��8>�p�a��l�����΋�����=83R/��4�c��Kg�~Ԟ
?���ct(w�:�+����x�Y*�����"���	�T_ث���Gk.���;S��RS�j��ͷ��ɴyB��_[����#�{��e�!��k��1f�9o��N2:��Ǝ���V���=�36�`WO���5�ӣLw^�A���0#�w_�䋦c������[7�����f-3�}&;z��� 漹���V_ ��%��}T�5��^�ug�	2��|�I�/(�| ��k�)4��П�ÿ�(Q���f)Z�40��v��]���i(�)�Ùd�q�ɻ�Q������E�+Ɉ|���x!�yR�w�5_���j��b��</r8"~	���2��Ɋ&|�O�9aُ~9oۓHN��F>�Qh+"���h�ph��_H����=��(�qs�G�Z�i<����t��$����䊝I������2�y8YeY7-�~����B����ڋ{N��?=�}dk���mu^�y
����ф��e,y�=Q0�y���*!��USF�����T1���A��I������i�j������Mb|x�RMH���l5x���*[�n<�&7�a�ug%��R��Si�'��������z�ŝ�F������`.RǼ��{-6��;W�Ō���F#�0ES���u���b��ퟣ�*�.�3\�\Ħ�=�PB���s�z"f�蝕�[���O�I�O��~=W֦Y��?W5O<��ru	8�H�#�P��?��8������(V�mv�c��׹0���\�{I=��� ���/ ���"�r�4͠�2�����;OD����0@(?��J���9��S�3l�G�Ms��%[ܟ�������g�5�~hp*ƺBU}Dɧl�0�4����tK��EY�z<��y�q�d�N��L+_�Se��fs��[=Ȕ���_03����R�'�eS�g't&!�t�al��H�ji�h�a�$oq����=�md��e<#c���D��B�I��ħ���P�}�h�1�"ן�]"?w�8���e������������9)E��K`z"�����#(:�J|�}#�Oׅ�Al��G�����I�K$�<t���j�I��7�Y:\��E��h�"%39�]#V������- �P��_�e%K���=�5e���2���P�Hi>�/���"=bi�*od�!��?��6'1o��kl�M�A�"��Z�LpB>om(���,�),��wN�.:�"�fa�]��w�`���nQH���m��$g�NӮuҢ�+_[=B�8�6�'<S5p]�KE%]��.U�LaH�ϤQRČ�'T8�W>چ~a�Җ�1Nǥ�"�֛����vt�8\qy++
2^"�]:N@��O[�pVz�<W�^w]�=�&�E̼;jzm��׻i
�����ؠ�񰠒��ɽ��n������b�X].M۵�^��>�+�N��:b��U�.![�8�:��|g��w)!�y�jr��H�a����|-5y��*O~�ݯ��[����n�K�(�����x�a��bP��dN�ɐ/�"mt�V�ޖ��
K����`��*S�������fk�#��1�{<H�'dT0�	d1o;��R�S~.�P.a	�D$Q�N�v����AT{t��~�vt0K������9y���gʼ�n͗�ev�w�8�uQ,�U����Le��I�bP���>e�����>�O�3�S[8��_�*r�ļ<�p����+��H�1j��t�jη�=���p��x���TjAQn���}���.7�����p�E�v��c���^�kI��t�Xu]nr�m�&�2tY
��SB	���<�qɾOr�w��?�c�J�2{��x���Fϥ��x�u�$�jv�-ŧ%��L %�t�N�r{4�1�L�t*���KX>����g ��ǲ�}��j;�K�CK�Ī���N���g �oYB���jZ-7)�2unF��1�zV��ݼ�Ƹ�N�ju"9��W�@^ᔶS��q�8��B�ȼ�5!�cJ�.߹�x�(Br(��ϋ�MI�b�hr���7@�E%����I�G@HK_�E�9���?s��X����-�7�4�0�d'Fh��k�(�j�����<���W ;�X��S�V� ��)�*tV#��dz2cɧkJ��4=��m��\PK��t$>��]{&�/|�C��dMA�d��V�x�>���ny��� ��i[����<"o_�G���w�0�cCNMTOK������oӷ�Z�O�S�׼$��v��$���S7U����ti�QKO(�� 5��]`P{,�
4���}{-�:�R��z��Cs�w�����ӣ����9=pK�Z�i���Ku[��;!�9h�-q��U��W[�r�ѽNSŎ�iP ��/�̸C��X�뾷���S�1�����,;��3ױ�Զ�s�FޝɍU�yt���Q�z����Z@J�&�ɬ祋Ǐa��x~�(j�~,����~�c�'���w;�"zޏž��juL��m���f������:yp��^�����Q���"��ږ��:��sJ�������	p��bp����@��>��V��Z+WS
�E�>�]����ϯp�$�m:�տ��U�Y.I��
H�89w��b��q���S�t�����"�qb�po{s�->��{i�8�+i������Ё̈�0��7�����L�-���i5��Ҫb܏���_2�ū��*2�ThѝJD�N.�N�>hJ낲Ҽ! "G���CGR�ZǤ��䢦LB@����!1�� �z2�ӭ��^@���;���X�����S:m櫶;p�b�Փ�{}y�I���P��F�p�����c������IWg��v3�e�F��? �y��&�޸OU~�y�=Җ��S�"�o��a�m����i&|�m��˝�J�_��]<����N)su��zc4����8�}�W�C���
�F�-ݽ�NG�7�m��j��K��A� �|��`Ϡʛ�3Iq��,�x<�0�1&V_�q�ܻ���=mc{X;�x���Y��φEY#8�w�sT�v�F���Si�0VS��t�M姼������	�����f� L8Ċߑ��|��Y�bb���2$W��/=�����2_v���`��$F�j]�s�N�p��ým��������P���H]�~ƽ�(�(���х���j��1I��>�J.�FIÆ`��8�����e
\��Ď��T͑<�htb�D��o���	i�JA�al�b/����&2��r�-!�����E�"�M�X��D�7�oW�ߡ��H#�-[�NN����1�n%ĉd�
�L`�X��8l�ȹ�>k{�����@-�:=�����I�5j��<��R�d��u"�]k>����#�w�f�ũ��v�υa�_�pl��G�u|���lcP�{� �-�2E"'���,����� ��U���=�6K�I��5�&$�GFR��DG����O$Y�꫖��~��WMv�?]�p�>h.8�E�l��%]	#�F�kg]�e^�E����q'i�y���p��j��:��U�t�(��c-�M�"��Z^4�0)�E-Y:�X��)o�I k�M����wj^>��'Ax��M	ʷݧ�S¿�k!4M+�����o٣�F|dc!�M�s��!�_L^f��k[���-���G�g{6:����&Ri��n����ΰ)`E���OCY�69����4z�P0ݳ�]�N]�h��҅8pI�J�iH�l۽]�Η�����\�ú7��T�v�Ƶl��#:��e��M������牯ٸG.m��{v.����zћ�!�1���
��a�y=#z���y��Q����],���ۼ:�:	�rK	�y��ڠJ�'��A�-m�;;+C�VF��K_r΀��`s��]�쾳oV6:t�+�1�+�E��/KΑ�->��t2.+m���v�;��:��w�)��T?0�y��W�^�Iu&�ʕP͸��s¦�?P��ꠘt��wɼ�����Č�F$�&E=4a��� J	�9��$�̭��u4R5�6�.}-����q��0Gu�9E��U�}���F��aҪ3��J�Zۛ�"���{�@�74T�0�Dl�9�qV]���/<�����Z�P�:�>��r�D'!�Q}�Z�x�Q�P�ꤠ�jf��eR[;ü�h6+3J6xj�7�}غS����A$�mT'�t�:M)|}p�N�,�G8�+A[�aL�����Fnв�+������wP2�5���1�a�x�G���r�\�Տ�vŻ�Z�ޢsj��L)���J1Q��N�B+gZK�h����B�*�%�w�\�j�4��Ntz`��t��;�։DIH���t�˗�G��.�ݿ�8Ig�h�\c���6��q[J��_�[��]�p!�?��|�T��#����Hr� .�w�#�#_xHA��7���T�p̬���5�
",�w���/��E�tV/~i_�%��C v��ne5���0�ʹ��:j`W���ޒK٩s�!�:g��dd?�`�T�5�9kQ�W�ʊ�Q-�� l%�S}��>�=��'����=�����G�(%�oex�K����!��:�U���������zH���yd_^�/\�(��{�M)^*@)��hw���?�I�sɘ(йy�kk�Q�m).eg�s^QV�l��@Ux�^��OaC~��֕�>s��o�n�T��T�%�y��qB��
��,�S���ۺ��vcN�_k����PT�	t��7���g`W���l���Dh�'��HI������_!��u�b�{0Y��}'��|_��O�J�����s%���N�eDh���ƫ�U2���Ϝ�!5+���\��3�9�է�P��e"����r�����}�$4V:�@�(k��漃�T��h�3�*;?=�_��j�G�Tpq��t�Z����2��'\��Cz�T+�4�>����!ɭ��7��Gv&,Z�2�c��[�
's_	��7���&"BK؈�J�����
~��We�މ�w~��a�L�^��G�L|����zGΏ��kx����`c��cؾ�+�i9;|���r?�`'����IF��A�k�>�fk�ʻO��Ə�G��DK4��r\��e<��(I��,���E4���,#�����p��X_ilG@V+$����� ��i���-nt��a[h��>C�Wv?����p9��0���f,u]tƆ�ә8�9뛘��ӊI�jO�a~q��e�#'��.�D��!g���!kO��n��s�0%�:9��!�r��G���wpӞ4>3nZAS�8�*�juS{!Ջ�0��f�^W�:��w���������t�9h_^\�iA�ۆ`��jSZ�7�݁ɂ���У�AB>��51,҉��sJ�����F]�<��t��q:q���W1ͨ�g��ө�
GB&`�H�!6 ��)�c�P�z[x)�ud|���!)ӗL�G���&��e���#��L��P�=i$?gnVz�k�g� �h�������@I��뿷yTr��ҍ������e�[r�N���1_B.1�-��D؜���6�鴎� ˵7��8��c�6�p{h���PdEevb)�c03�-���Ɇ�0����;��ҷ�z�{�#:�(�^�ud���7x��0����ΰ�f)	-�?b�e���2�A����lDXD��BjIǪ�=X^�e����ܩ��/^/OUC5c�ΕO:�Z}^�Antěa�a.i6(�<��ڙ|$K�}IB�(������=�/�ͯ5���U^T&��Pb�bq�'��F�$K����.�IC�9֌��#�1w'��۪�^��h�g�]���6��⛆QQ�3��9�u��4!��;�b�(}_L�dJ;��|;y8~���-�IД�XԖP�鐭���w��f�?�m+��!���7s�:�uC�m4��|��V�˯�?py@�S�q�_��?E#��W �s����M��P������O�2� �a�8u<������M �/Z~(#�9�!_OCo��������r�BSb����-��\ߡ.V�T�f��etQ>Q����J#Q����AX��%��c�!����(8�������'7:w��\��J1t��+�?L͢�z>�����	�"G��.��\w>F}��	�]l����=�S��o��~��p�e���	���/�J@x��T6��T�����7.G�G~v��j���g)�c���0P3_B������OZ�X�X�kL�bz*ͅ�����Y�:�5+JqDR�a�Ms�:�Z�(���+��.�m�|�r�e���梌~�)��u,���)=�!滅�[����P0BB�CT���0�@Iw�R�)�ٸo��z1^A�{ch!�Qy-ݚ�ɿ��t�W��	���Ȳ�k8��PM>n� ����n%��_�7'�C�yZ�v��a*��-c��GB���ES��[-5���'�5y|�n�e��C5�1*�C*e� ���	��`��PjJ�\�E������'�\��=�wԆЛ�!����C��Db������Fn�i�����ʣO�hm�K#)D�O;����cI��ME�Y�喖�����S"�u�:�ը��a��<9l	�4|���/�e�� .ް#H�X�����p��	oX�1Qg����Vz��`Qi�I��.K����L7�"��|g�Gi�g3({���p$�"�;؍��� ���x����O��;��K����:/Q��J�@����"�ϼP��Y���_�Ux��_�B�?�q��<�MB�}�o���{��Y��d�ԧ�p=�x�a�߆(��㐕���b]mW�gwAn(��Pohe羭�9EZ
��k�9���ޫ<��O�{��mE#���׼�PrH�&��g�V�K��dI�R=#��W�b?�5�&�(�GRZ��fYZ6��?��-ПWV���c�Tõ�0&�6ߏ�u�`-��A6�#%�� ʔe��i��ӻ��/�7�=���ŭ��3�G�~���Ȗu������#�w�I\��й��!������o|��;��:;���3��}��)�D�q������k��u�k^e����X�y���6����XW�뮇�>�$.@:�՘Řn�r�nR'�I�Z66���[j�'2��@�,�.���nHr�,>�|���B�$ v�	�%ï]�� b�N՘��`��T����Т�*ڢ�b�Q��y��р�xS�.���H�PB��ɓu[,�nנ���~�I��'#�="s�g�n��Ѱk� �:��Ӡ,�"���!��JJ�3Լ��,��/'�<�\�,���\�H����m��a�'�_�F�%s���
�
�A�D��n7�X��Q0��6��2J�^����|x
�ĸ�� a��y	$��ee.���RB��������4tp��گ�ash"!��}�	��$C<�g�v@��9&�:��+�9�D�o��}��/��c�$�Zw�8���?����Y�L�����L���tR�@���	pT��K�ߊו�gw6�w!X����@
�Bs
��OK��g$�r�<Ri�T.Rq :~�91��5$�U�i���QHW�m�4n��L���w�h���g �_= *���z�Jc��ԛ�N�C��=���|���< �uC0�d��`����M�F3x,��y��VѳE��ݜ� ֩8�"&��8�3���9֗�R�茅�2�3�jTS��/�N�ݯ�\��6�#�趔T�`�@p��=�$T��[��>����_:����pv����13�%:�2U�'c<'�~�ëݧ���pmB��� �=*�_�e4��L���ImP�bµ����7!�
�O ���e�3��dD�cV�yU`�������[G�<�*x�"fޱo��i���м ��U�Щ^��R���`�����l'�V��H������}�q���L��k1n�9'�>g��9�k�L[��`"B���C�e?N8�YR^H��>f�G̲�t��+��"-�s^�Es_:��1��ꎿ�{v�8�}�p¦�+`��WnX@��\�����Hi#9%8WWG���x
R��3�8�i�ug���ܜ���T�I��3�����/�Y#�����R�!�|�M���~��&�3��Kv��	��\t�t2��I�����t��d�H#L�¾��m�,== Af<!P������~���5d#ߤOF*.�Ó�5�	��wG��n73Zn��D�:���Ti8K��Lj�$-<H"!Ѧ������n�V�L/�fr��O�6�OE�!���|�M�j�B���@־yy� P7A��a4���[m?h�Jȋ�:f3�C��#,L������WP�P AR��<��s���ⅇ���/m�=O_�F���gY2�����pR01���ԯ-x�̿�s���~�-ĸ|��]Ȫڻ,D�!8���=�'�z�%j��r~�kR�[���%~�i�$���W�A�x
�w���$a�ŵbt�"�Z��N�������+�rXnV�|	�v� ���S��e����嗍K�Q=V�yr&���?��!�� y(�����J��ˋ�'�������U��<��1�
����>�R&���r�����7�O&����������(+��̈�Г�}fr����'ﶺ����g�v��<��"
~�h$F�:p��+�MԌu��R��%Ni2,_�"�_��G�#g�D?��P�����"E	��cZ�P��$�7C⼬�15���/_5���J�����B�=,�ѧ���_�؊A;��B��2[�`��;����]٥+�
�o?4��5�c����Pf2�I�_����4�b��N<����$��K\�ډ��a�5��~U�4�:0>��Y8�������kښ��)�,>6VK`���r��଼�� �e��15���(VH�s���I��TɈ�����E��ݶn�#�.�-7�c͔Y�n��� Q���?:��T!IC�z?[��a�b�\�z�/]�-V*4�؁؊��h �j�3/L������_�4L3�Si똎q�rIP�λ����Ó��\q.[�1s��l�Ӽ��Sd���ۻ4%�\�T�t�+ߍt8d�=���w'�h8�x�(���"@�O*7N����;�2L��B=gH�D�?�m�8���e��(�jtt^GC���Z��I!�v����mS46��O�
�������&��
9�j[���$�w��5��!��h5�� ��
Z^�al��.c����A� ��ˏ�u����V��r_�> �lԨ�MY��Q����*�C�}�Brz���1DG��� ��Hu�Bw��> [��=^.*��5+~�#u�&�ng�.��2P\�j_�f�t�zb�$�q�ON�����>#��c�]�Y��@��5 ��.ARtV; �s���2髋�/ۡZ߇�����Zbo��?���>ۼ���l�A��~ְv-���)��T2 z��v%XC�JpT���jE���@�$�M�x�Hէ����1����<x��P�f�zk|���`���0
@�au��e����ْ}O�hw%�Q�35�w��d/VC%��
MӶ�VpXI��T�c<O_9_�D��	�z��&�[;���a�Bxq�:}�Z+{���Y�W~���Gw�M8(�뾥�<NC�Y����<Q�)��JB�=8� �L�)���	D�	=���-ޭ�����&�V�S�P��+��q��H��A�2������?{�e$,��F��!���e�(��}�o���{���ॕ�~>��v �9�/�v��o4�kΟ�s���G4w�/Gd�s����_Lvyh	�}w���1�M1N�Uߣ��ⵛ���Dd�N����:IE��t����܃��ʵ
���~
��C�^Ay~�[�?G�����g��#Z�Ql�<s�E?d!��>�Fk�s`
"G�S����5���3�T�Z��7&y'��x� �e��{	x�Rl�[��<�h|4i����0�W��<�x��P���iiIk�S�pߜ�e�Wyb��`���L?�b���Y�a9�K�����`
$zMr�U�7X�4��0K{s�5Wl	��n��XD֡�'|��v�ߵ�۠3�
�B$��>	���.^gk"���H��b���'�<!��'lQSk�=�Ջ;��	 Z��	~Ά�x?b
��8���J���R�;�Q�0^A����[z�{��݉�g�V��QY�e*����y_�l�.G�bF�\��Si7Y�[���&	��J�����^��6Ɖ�ot|Д��V�G�;�Xjb���#�~I�}ٕR4��I��1ѩAF��N��W��B
�k_0@�T�dKQA�� ��w�~Xs�s��3�xg�I��a�*��m9U�׽�`�����V�ʝ	�*9`� ��� 2��*�0xN� �u>7��U�j91�Y>�D,��i9�����ݏBU��X�3�ʃ� ��I�-��J.��"Q�pbl��mVBn;��TlZ��2ej�Ѐ�;�/�X؅p
����͐�_ɡp���ʱ�R��Dh�� G�<�,)8�=S�����J �تZ�j����X�SԸ����z���\���|fL�����:܁�qH̑�{�[=[,��cA ��]����2.W�\�j��q�-$=����"� ���Ŭ�V�W��:��uà'�ۗy��o}�g�pȧ��}ͰZi� K|���A����;�3U�}�/'r�냁�fU��b�gT�i� �B���*@V���L�ӆ�|�/N:gy��ˇ� Y�#�$�Q���/I��+
���wz�:�sR�6�o���<���	�dt�6�}9�]#�d��	��o����-K �22}�Ӟ�e_��eLl��Né��2B `^|�ړ6�V�(�c��-�4��t6�~l�_kqP9���3� �RKy�bF�1��Ԯ����w0Q�>]J�}�HQ�����>uS{� SF�ܩ�<A+z��o?��E5����r��DX|�������9<}����F4�mh+�xyU�<��>]���L�o���|T���;\���x�>9?1�>$$Ç�{y�������_yc���`�.������x1����pH�WMZtQ@��-�Ñ��iY1-�}Ag��U�@�n$���I�K��=��(U��/�*��0����E�߻�h��ޕ�E���������+9I榨��le H[Cb�^"@�AU��v�/�8B��B��;�f�/9�CA,�z���=��"E�w�2��YҼ.:�sY&�e��13���⃱ſ���Mj�Po;�}elgrM����`h�������J��9},�n3"�����=���W����ʨ1��7�M���ѷD4�t����w�r�X���Xl���<Ts��^2�� f}􏿄��R������~ ���ԥ��2Øi?Q��U@8���l�Y�o�����¥�蓼$��%V ��z�  � ��zY~�nGU�z��W)��$3��;-`�U��Oe���w_�)��ȓ)�~Ѕӗ3'�%dg�����V���Q��z=�&�,�\�ֶ6��KӇ@��I8����Z��;Zd@b��y�4�dνl��ɴ�ه�4HCM��=��4 ظ߮�K~]q�9P]z �L�xm)��-�-$��{�=�̊W<]ꖮP��'�֤N�
 �eh���iqW6����4q`-�����H�or��@N岥��?yJ�T��HLo�Dш�,d��(�G���F �Mom{���)�~��E��oԏo{>�tɔe�)4�y<�h{�n��${�B �	P�\�Yz6&�BB�����0��	�=�i�Y�^Z�^����}c}����t������+�{_�,F��o`D�'�� �W�]U�j΂�������_�Φ�go�V)5�M�N�|�"�ad�&Q�(��'w�GwhI2A�.��8f ^�J����|,�{W��w��J�D��zq씂��n�؈?9�x��� ��w|��P@��ޘ���}�px���c"s�L���e��Vi�����o[,&�������U?��'�Ȏ�@?#�w�iQ�t��Jz�A&�8�5�՝�m�w�<o���w�f�P�����n���R�U�7�KA����;?Ȣ� ����Zн;	��}W%��������ؠ*a�ѧ+�����x�i|� ����p�j^�2��kKZ����Uc<0a�L�p��TpA��_�X��=��rи��ć	���9$$ak5M�v��GS	��k�%T˶��?Z�n�`a��[�u����Jv��� -g���%'|U��u������Y��^�ߴ]�|�2?\�7Ѓʘ�3�$�7�����9a� (��6�S�y��Py����	0)�Ou|'@h�����_��6�2�F��9>�_<��i�Z�Y�u%�?�2π
^e�J,���' �N��om�n���N�^�F<{!�"q����d=�NwߞOm]d:^1�P�ޠF{�d߂�9�aMR�?��C�#�zv����3��iO�ӥ��89ٽ8J�!Uw�,�� ��C�2uk��y��>�qC�7��G4UUbK`�Yw��$�PL�i�6[2�}:��tg��H牙jcv^���+^�ʐ��������]\�x���{�mO�^Kb�?��)~5���p���k�L%��m�[@ӴGDG�vv�t[}ʘ�����*��<\o ������wu?n���3�����|����H�3��/є"�:�ЏpJ}%B��U���gE���A�-Q%�BF2j<sX�����SIL����\�C������ꅔu���K�r(���3{S�ka��[
h�=�ۼl�;�6[S�{��w�[�0�j ����!>���|x��ǅ�,aB�f.��� q�����o�������f�3�yp"�����>� ����Z&_�<}�纳�壄�
��i<e٤��X������k�s W��3�_��-G7�aM2�t���T��/҉i3�OZk<���Ѳ���<�`3�����'n�5��
v��Z�����ۄH�_�X�? �=-8zg�v�hqo=�B[,�~�M�\},��z����s ��}��C��Lp�7N9��S�]�V hO�<V�1�!����!3?�zD�,�VR�=�wcN5�SQ�P�'���p��|�;�/��t�q���L$�_�ks�^����T��� �t���'t���..�W�G�@dܞ,��6i�J����lm���A�����q��ɀT�id�e���G"�[����8�u3Ev@��K��T��6[�)�<s�6�JT<�A�p��| lր�8��LeM��qT��#�(�$�4�E�%=�� ~	i|9���v��Cv�p�jb��tjP�&acJ��D�"�`,��b�I٫���Q!:ݢ����
���<��4 ��w:�?QR R�Γ��'b���q����Z�L�U��)�3�N�-k��̓��Z���[�
�����O����9:@��6����_0@vp��\'9�Ѡi��7�=���+^�m>�h��2qx�����W�xY�E���C,��%+1��V].3ѣtě7B�BG�&w���?E��!�v������זl��&��U�
π�5�'��~��� ��F��僘�@c/���JY>�)� ���@�uK�����<��(�)j7
끨Q7��T9��B*Ap��&�9'\�YZ���3�c<#P[�O���o!��P�m�~�>�O3�����h+f�P�CѦ<������� u!�:եj���>�M� E��n>E{��(�ОE���X�I�UYَ
R��d�Jjٮ����a��+v����<t�	��� ����]�z���zbI�F �H����ˊ�9K.���V�Ե�[t��9�({h�����(M�ō�X9���r("�mǻx����n��{���$��Sό��O �Ώ�@m���MHO��2%:��!	֗Q!&���1��7Z�F/!/d���P�kOz�SB�|͡x�I a�g�KE���I��o�셇�b�i\�Ep>]:x��V�t��ay����(�}�~s�ȱ�鏇���{h=�'�,net�'dZ�4s�"����n��T��/h�Z�j~�rD���H���a�[�)W���s�[��0:���4rb�ʳ"x��aQ���@�Ĝ�tMAf���ă�W\R�������J9��ap5i��fd$=q|G���ˡ�	�~bpr@��wm���M�K2�6۞ylI[:�vk�^(�n��z��mC���r���-�T�e~ӕF�K{�k��r�`e�=���������t](���(K��P7%������S*���No�"$e M�ˣR����u����F��f�<�\��v��8��L���>! �<ȥ�|�f~"!��a85�w�m��7x�^��囝��G'.�ȧE�<.�P�z�&����SyS���z�CX-i��Y�*�A˾'Pf�Gy@�>���wh�^�3��f,��f����V&�U�U	�u��v�b��[I���ǜ��p��p%�����7%���!`f�@�z��㐏�Q�UG忲��$�}?�݉��8�}�kb0���'��@���*��(	}�/7���U8I#LX��hC����k�~��\}��'���|�Z�6������;O��κ��MivޝS��|qq��c6�\�G"o|`-�[$?��Ju��2+,�G����[j�2�?����*Yu�)�����k��e"�OzU�#��yJ��bh��v�T���x���H��oi�fOQ��^������h����7L,����͈���[?δ#J��ֵXn<��l�0�;[$������'�)�ߟ�38R!�ۮ�^J��J��5q�d��~<�
�ʈ���� HxSLY���cl� er�3AY9yE3}��	�b�2����D/����5"�Q�7<��j:UmwM���9ڵ:&>�!>���J�ˮ��-ޘ�o9U�J}G7o�:F�B2�=�Q}z-�y^fO��Sx��ӷ�V̋����ķ;r{�����sz=�V.A$�-I99Y�A�o��d+t)�D�B���!ql&��l�2���>)�4~��e�.ߧ��<'�2�@���~@��ՋR)�J%_�m���zT�4p�{�Na
�g�mh�,o �\X6�1V�����G�,B��_U6FO|��-�8_w�9���.�5�5���u����z����v��;��������h���D��/�=�kVb)�^�ߪ�y�,���P�|��ⱱ`L����O`f���;-���53��~͙ަ�1_'��L�\z�٘r��3�?�_��m���������j�c�����h�!.S٨=1�q�H�~v��������=�46�U�V�}̽t;�qc���s�X������_��O��O��Or�o�B(I��i��sXΟ1(u��+`�;Ň1A�琶W�LVzB��t+D6r���ɇ�Ҝ��;�*�aw&����`J��NJ^�б�
�1�dG�v���13��]�ݭ;���!���e��7p�NB	x+$�F�[��˄r��M;��j7K��ϋ��@nM�S���i���JgKL��L�\�G�t4/?��I���:~٥��gN&h�ڣ�a���#�;a!n)x�I�ו[���K�<��'F8 <s�΂��G:"���jY�3Fܬ��/�J��O�*�J�!AJ��i���w��r��f�ݩ�	��[�R��>�|��qﵶ̳�&`��ZnM(��.j;%��=Ҁ�1 ?��n7g�
��˘؛ԩ�����%'D1�����}�����D���Yf����-Zn�U����v����+DQ��w�y�"�"z��<�L�oJ���qZ|�75�;r����k�+�����T����V��[�o<Z��ɫ)N�1S4��G��E�c2���������E�N��+Vh2�s�TH�\k�����5ؐyq��U�?Q�:�c!��O��~�z����Q��82��^�
�пSBW׹���n��g(Kb��:>�#�����6�Z(�O�mk���\IV�5m��KO�"p��PɌ|��>��7Ύ�ɚոHh$ҏ�I�\�4t�e�թ܋�ecIʧl3�vs䘭�-ҏ����N)S�q���C�S|�ʢ����5�l2e ��� �	���f�r�,�����YG��<5�,�:uk�R�V���*���y�0`9�ٖ|56�<F�� �A������*�&����^�]?x�͚��s�b�7��O�Q�
�E���{�������m���I�!t-@�����ˑ�E�.��n��h���%�����H����9��r��//8Zz�TYr��V~��?��_�� �*�uȬ'JI�)7b�衮 q�������e�tO܁��oA�y���_�V����[�����|�8� ��Y��#I[i�28�K��<�����#2@94ܾ�1��d�}�^*'y�Z�TH������,�1�����~7���A^^�
�E��_y�	��Gc"��;�����Su&0�Gl��I�7�=����&�Q/�����"�}��޼.*�����BIB�a��97�����r��`1/��g
_z�Qx�4@�g��搵�H�!�R�kg>�3��lOD��x ��v���WP���I(�����jya0���ฉ��B/i��.T���4�G߿VT:P�*�<�R�R,̫�|�Dsؔ�����:�aK��M������+F��`�+��Y�H����E�A�z����Y�'����f�b�Z��*Bˑaռ�ʪ�?,~W���mK��S���#��;��bbh���( ����9��l�h���/k6�}��#�'S�G6�n�֡��zA���P[�}�1���g�����Y�4>�nQq�|u���ܫ����{1|��-����:��Q�@Qw�� "(�]�J���R�%(�-"Ұtw�H,(�H�t����������>�w�u�qv���s>q��]� u؄�M��Bw�m���Y<k��W����3H^K�?���p�
��G��ꫩ�VW�%1̢$I�����mC�����~���PD#�4�Z<��l��5_M}q��5vM/?�y����Ym+���Ӻh�&C�z5�-b��V�=��L�񰅭A�* D��{�􌔌�c�y���*y:��hȅ�uaI�tX�8�1��^�|(�Dԓ
�K^D�{��J+��U?��>��-��A���o��c2�qq]^-x�o��Y@{��rR(V�>�R�0nKj~W��pu�[ma*�W���2����Ų`8�5���!��?��l���[����/��O����� x�T���A��h�ϗ��� �B<3�c�y��s����;��E��r�ҫ��3O�~T��Nj�E��hJ��L'��W�>48-�GB�y~s�����o�S ��E6]�.��nk����w�_  ��W{����I�<�g�D���bܡ�h6�*���G�>�˱~�M��ydg�iʭ;�¡Κ�g���A� ؊g1t��V����(�g����dS��4G���l@�4��/yEmd�^@��]T�* ����+�fm�i��K�u��Dfg��&v�'oE�D]FQ�l:��m�(
"X�g}��Z~k���FD�ħ��P̚�l��&���3��4���t�d�D��8����2~�y6�C6�Nfi.�7c��� i�8�СE��l�������|���/��� @��"4~V���/�_����:�:���2��$6� E���g@�lq@PA���\��j�ʮ��1��xƏB"+��[!�@�S��Tۖ傍hw�:)˗4�5!�C3��FМ�*v���_�����N�-����Oo����k�'|�
��nŐ'q�A��+����8����n(&��fϘ����e� ��ۍ,� ���ac�"�s��9
�<�{��In��>9�	"����"��Mt��D��	��r[#�����ڂ$��դ��������b�P��AK�V	��i�q��`/Ɛ�2���.z�����������Y�Z��\2;ƥv{��ܺ+4��L�Q~M7KȩK�f-�~��&�	t�o|�%����`��E'� (C�٪�LJ��gy��pq�7��O�ǿⴿF(����4��?+�Uգ=~���֣$a�� �n���@P©ϒ����O����9�e��gˉi�z
�U|�mھ�h��eй�dN�E+�������Z. ��秅�ƸČP�D�q�il=���Z��v�a��PG�!8�32ܟ��A�	'j�K�|�˭��ϳ���I����/[����8K8˳�ᘘ<)�V593N궷�a����q�}}���+�o-m����`�ot#l�b��YgP胋��p�0��]�+�$,H���J�f֤�qH ���������GL���$�:"�0�}���C���?��I����5�[��m��" ɶ�6�Z�>p�D*�aqJ?|vȒ�ߵK�pt�݆��
�E�5x�E'��R^�9<c߃B���'�.�7낔�f�% ���C����̇�����7�dr�����Znt�	�T��a�Y�F>��E�p��vǎ�_m�W	���^i����	��\��f\U���tJG&f��"������J*>�9x��\��nRQ���k��<��U�����/e�*�/����oUޤ�hŧ�E]}��FT �0=;�\jE�o��'��7�-������V�e8���X�"� H��7o�y��}'�65�hq@Ő�Į�A�|o�R��E�p3�Q����X���r} ��{��������B�Ъ`�c��{_ʖs��vf�ټ_�xV�s'�� O��?�����;������+��_�x=���-�;-�&�O�ƨ�!BD�qnYP�w��T[7U+�5��=+ؽ���n
�5vu�ۢn!z2p+���:���]�O��������(9f�4�E<�W,�.d�>ϫ�)K�5x̭�Ƴz�R��Q&�3C�%ǌxS8K��#-&��u\J&�wu����ͳM��	��*�ć��=A��bI��o˅�6�!6`�:�<�~!�/�?�nS^�q�z��8nN�TB�)G�kL��2i����"�t�Γ")l<�H��cV׽�H�L�z)g����6)������$͌O�6��z�3R#"�"��9�y��wg��lP�dpֱb�����#�8p��)�c|Z�Lփ��P����D�@�4�Y�ѸͰ��{ZW��t5��Y���i���(UȌܗL$�'%��[��Q����9�����(���1[7��mPo-�N�$,����|��)�v7*$x.�����I?��3���_��䨗 2=^<m׿+��	~ʹy��F�,� ���ӧ�x�wA��`��:
��t��"�!�����[��-@~fA�Og�9虂Sg�fN�T*�tC��;%D%P��b=vg��z`�'A�uLnaY�
W�1�#�*�~ȫ*��k�h�f���6-ȴ62Xh����5��G����	֜u?�ʽ��? �)<30sn/�b�)!j(���u�׵^�LI��5��>?�8�q�K(�a9���Pm����Vg)���c�Ą���a��&E���~;z��L��p�Υ�%f���â�6[�c���8�����h*@��+
�Wiu�P	Iɇ��ݨ�^���$�݄��z�?�,٪B��6���X_�0r�6�Gy�k	��!F���G���Y��ر���5����Y����V+/�XÙl�V).L��h�����GHL�f> 2��r����@DK��i�����&LPS9ţ�������$��8�sI\�12e��p6I�����e!'������?�]��#;�?�E�2f;?��.��}:W�������-��DS���i�/��X�ƹ�N��h1��H>;3=�,6�FCl�z&�wxa8��ӌ@ek��<>ٍP�<���ۧ�4s/!�Y��|���%�.sfd��n�{3��>�)�'n��V�Nkqt����D�@��2hk��� YG�P:0�8(OiW���t>%�{��+JcE��@}������@7��H/
ݕ��+g��/`�%��ė��ex�C�J��� \	ܱ���"�l�Uc��zk�Y�b4(�W�:�;���^j�K���G��:@�Y���4�=��wK��;;e;kS��_i���ȴ���z�Gx�����tw��G�^t����Ond{�љ�W�A���益�ln��ɛ8�h3{?��Gu��Z�7Qע^xz|`X/�ƪW��oج0�����r�	�+�@����ʦ�B �3S��M�|̻�)�@�z��V��l6���=p�
�UC�@���z6��f��s�&p{�Z0�����5t��}�o��J^���\O�s�r���&Չ`�
1��M�a��I���K8��-����,.��_�������y3�+
�o����'b�a,�����T3Gq�w]�D��b"��*`��\)����?�yy���Wd�����
^J�Ӽ��q��/���J�3��$��y�����V��Ё0���_�N������We����/E�\�v3-�*�@�p��W��	�q�*��� 
-(f���v�z���LO�� �Weuw*�4����;E�@F1�:���Ŋ��!z�F����j$��sXk�qyA»��xɘ��S�)[���t�4�fu��?ɂ�C����cv.�{�m�K�4���`�S'`��"�IłZ�_R���*����-�Q�eb��(�?Q���k����SR�Uo.�P�����h�f��Q
�R�����L/����|m�a?�P�a�o�o'�����`�t��l�s��6��0��A�nQ�ł�K�+��B�o
�R� .FT�U��_�������~p�2�^D��G�7�� nM׫��\kʙ�u�v�V��=,y�L4Q��c�P��^e>/�/Џ�1rTC��^��$.��7�B��&DzYbk�́�Ke�s���r�ϡ��1֮88�^����Z�0�/����9ب�:�f"1��C;�@Y��d�B�}�k�?�9��������;��D&�Es�#�윂��U%6���!|��W�J��Ex_�ߵV���W�JMp�U����ݡ��<�5)�]I��NB��Ꟊ&�/6�|�x�"��R(��66d	�i�ǔ�y(N�.�����mI<�� ]�l�Y��T���
�^���]&�!o�^�H�1x��;H��&3��0�D,G��:ug4�q�
�$rM����#��{�0H� ,TC��iK�;�:�p���"��� 6��<��G2�i�w3G���p�l�t�|����Nv��p�����2<��Wm�!8�iH��4rN��L����!M�Y�r��e~w��K��`-)�)�I��J��Y�TH�j�]>D3d�S@\Y���!��|	aM��t3��O.���G�QgW���1���C�Oy]Ϭ7Ͱ/T �W?W�<jhG~J�{J�ߌ�TE�E�����AŒ�^/Z�D:��
���k���d�߿�9j�� �Q%А���^ܾ�.@Iz3NY8ш�a��SW����yǯ�gq
���������.n��<Rʇ��G��� ��V�lD}8���J19h���?O|Q��:�/�!����άVKH�n����c��a�Q�>�ʬ\�X�I5)-����:����;�;q�Dz�dgd�\�Y��wۀS�g7è���uc�g�o����4�k��o�b.T��B�$���d��o7�K7��aV�%�԰f-%�=��?ح�]XE�y���(u,��2&�+����jM���Q���K�����|��[*��\���8�� .XR�~��]���b�=y��Y	���� ��=��zkZ)�h�(sq{7�����Ku���ޘ��vl�T ����z=&9���>d���lB���o8��+z���� G�
�S������D|���"�:�C�e�74�Ɯ��j���D��4N"�R4i��y��p߮���M��G�n��*��
�/���D↭ޱ�Jca��eey8r���о24m�gi��ȍ��yѝK>�sz��.�0�iWQ*n�Y�i%��D�9�Ky'4�s0�8�&��in�w̧��#?����%�9�?O��b��`����6&�hc�Ÿ���|W�;�$G�'q<�J!]�6((
�������/N�u�ng5.�҉b�b(���J;4��2?_暆�+��5w�l+��t3#��J;�$i�N.5=T|��!����1�fD��i��� GR*��j�j!�]W��1HG3# ҕl���B�l�Z�Ǹ�}�5܅x�iL74�c~����C��-u���J�~݅]��m�1<_��1�X?Vv��,j���q�� &�W����C⣶�������X�/M�󯌝�3�73�1��M��`)�3i�WɄcF��>�]=�U�#��BY�D#�]ݿ灤<�8�:��S�� ��ǋ����9�ˑ8�;�����U/���;x1�*1��u���Z�V��PN(4��l��eJ)���@X��a�!;�<"%��<��[�1UK�Θ^k� l.�q�6�l��`j�%�K?����|��#%�|�P�43����?6%��:��e;�;�q./��;(8j���I�B���H ��gOQڔ0 �}�0l���J��͉�)5�ZM(du�Oê��b3�T�8$;�����+�}Or���o�a�a���߇gi,�]��O��?r����e��q.��g������+���y}�/��L�8\<�T9���K���|���U�;�Y���w�����ĀM"	�+�-�1A�3U�j,�jу�́���KNB�Nܺ�i3�n5���<<�#FZ ���c��3��j����f!0o�$ txF�a�Qх��������j9����d�c�N�\$�x2����_���u�ڤ����3_���PG"3�Uv"���̂��-�գu��pm/��ـ�_n�����
�����>��BNu�,*+�e�t�R���6 �<=-��^<��ƌP��M4�5��3	Jt8C"ud�}wH���W�!J6�/����H:��
�v�$�7s9~O��Rb��2��W����n�#6���5�G��Ks,���|6�|�5.$|�@PS� \!��?55�{j�XѲڸ�n��GzKP�۴����5�IA}�B_�Q��&빏G�Jw3�i� �\��~��]�8c.Ҳ�M���x�#����BKԛN�@��M�s���Th�2�v-�>M�*��Q�̓.�����4�	3TV3 A%m�a�v2G���A�k�I��U�g4"�����msw%qyq3"n�n9R�	��Ѣ���t�H���Ђ��l!�2S�T���X�e�@��Ć��Kʤ�h�*�p��e&Jy�(�Z2��x��$;������o5����4���=&��H駊�O�����g��:����V��874${��c��z�� ?m%P�n�?����8�LjE�M���r偦��].�O��t�tY�Y�|,`f�<�Tˏ�RM���H��d�ݘ���=򱥹t�^�<�IBb|��	|A��%�`��pj�(3�Ѫ����慖��w�r�	�!T�'K=������nV����l�O���s�3 ���"��u�=KL���qB�f�LJ�	
��5���g�[���/��ȵQ䣍]t2�����̻�/k��@��,NW%T���q@v��#B�+�1��jE|<��ҁ����Om]|�!R?*�hRC�	�zd���x۬��L �ʽ(AM4uu���'��&��$�2��� 'r4TW}II���5� ���xB�ߩ�������yJ�rJG�ԟ\�}:�[�*.��GS�m2����O��H��?ؽ��0�~+r��GU�����"OjC�i:�$y�3�a��߱^T��2��X���u-$|fd��&�KT�1�@F�N ZYٍ��A&���9e_2�)��\�@�'P�m3�].��1Nυ�2��P3��=�$�F{W~�a��
C!yg�u~���l�FA�JE酏TK�8���!]����eXcW�xxn`u����F�5C�C��D[�Q�pda5��5��W�2�l��޷���_8)]MV1g���|ȯJ[~D���N�����.��7����@*���]]1�̔�%\��%!��������lK�{�KP�ɷ�ٺc.��7�Iv��9��IϪ�?��7V����+1��$b��HG^E�A�/`qdN&F|ϙ�Њ��1�<�*��8��&7&�` �Q���p)�J��\i�w��r�cŰ����.���<�B��7IG�h.���b,�b�a1��-.]�����7�@X&�jb������DLPf;(&�lX�%m<N�p�,��4Hx��:Q���gH�I ���(Y�ٔܚ�>�{��2S�=��\Y#ݽ��O*<̯_p�V�-��'Կ�d빃�(5�MdWV�m0Nu��RF.բ푔�� ����� $Mz�'�i�L|���R懇 _ͷnNGQB2�By���_�7^��6�B���rrX�B�r].�8�?�x����C������-�3�{��Fk,�sI�,ޝ��D��i��D�L�M<Z��yM�L|����Y�!Q������� ���L�H_����yR�%=����:��z8n.�`��s��)>�@������xV�E B �V'�ah�)�j~f�@X5�b���/�k��Xu�0?�r�����J�nM�_�H�=3�;o��ž+��?��[��0_��т�O�k�^��@�+��fՊ�
Vj\X>V:��:�����I_y�����o6��\��A���7'2//s��mA�k[�b�����9�aBX�����5�s9�!"ƂȘ�6��f��p�s�Y3Li�D%{&�����I+pAj�nݮ���C&J�p����&��>���9��G>p���;|ֹ��-r짿 ��<�y
����gCX�-���W�����Y��B�����0$��!-oT|9,��+�Wˣ����k� Vy�w�H�Aȶ��h%�j��?���{�B�5x�QJ
^I��,xވzt�����|�I�X��7���-�d̴^�%ngCu���Ě�S�����i_��s�.�i5�ЀX����ĕ�s�g/ �F��߶�U_�rƙO��������w�	�5��<�q՛����<�D8E,V��Ǧd�S��{��YXl<aRh�����5I�^���K�f�`�ֳ���3�2W��.�?���8��_+P�1������M��f1j��B�?�UH��4����� s��S�~^���K4��=��Ѯ�1c�3��L���)���K����e�Aa���g��qZ�Ti��_�����̷)���������E��<�ȭ�K�2n�)��dĴ� _tUQ�� ����r�?���xh+��A5C��N���K�.���w|�����3�IM��^t|�F�^��WSs�q�홭����6q�i� ��Ĩ����N��sH�=��P�rD�h�����A h�2 �OӭgJ�d�MH>���j��e�Z"x���hz ��;DL����֚BC7�Y�9>���g%A��ͅf���:`'��p�\��9"
�E�]ic%K���j7�$j����Y�P�!���t��؟
�
��X-rA�o"��e <U��SHu+4�¼|�m��������n�ɣ�2���N �G��wT;����d6ku��uh9ܟ�WT�nv����L��� 
�L�u�8�U�E%Iv��||�iS�* ��E"v����v�6��j������R���; U���ܶ�pb�I� F(�����d�C�,g>�5���wݞ�,�8u~�>w�#":��L�b�Y$Ԥ<d8i�q$*D_�����h���M����1౛ICx��g^U��Q�,��8 ���̀�p��mg{|s�2��Yp �J	P�:���s_�E8��N��? ���a��0����e�4H�cz���a;~\�ϻmu�A���ݒ�g�1;P�K��B]K�͇[���՗�{���M�<{Hq3Xa�ۓ$7>���aTh��	߳3߂;�1?��٘ 
n��@4�6f��  �ө�	�������i�U�d6�M{��NMK%�}5���)ݯ�.uRk|U��yj1�j���-������˾mA��G%>d��`��k\��Bo�WY��)�9�y��fi��=��!���a5ː�?6��%u��n3��|��rf�����t�@�x�FF4�69�1�x�D�?���,��6�d3_Tl�*k5�m�g+�w}�\���K����j-��[M���{B)���M�L�V�L6���;��DP1%n�W�'� ����x��" =q�q�p�p�����B�c*z��'+:��Ϝ�d��&�;�:/=�tCI�1�I[�D��رw`E�>i�:��A Agz�K&&,���1�,99��)k�k�6�ӝF�v�Q�6<6����|��P�4td޷^�i1�Z��"`��r�ןػ�2�Ñ�8Br_B�⏷�)����T�S�X�{|�y+��zgL{�KƶE�>~�' |�65�����݋�b�����D��i�45)II�����4@a4�6���1C��#�Q�ҧ}�l�G!C��!9*�*�b#��cZM�mZ7�z�[���
.�b&������ D�#��-�\ڎF1:C�|*�P��:�x>��)�9o

���ih�����^-9"O�]Y�,Ii�'@)�W�8m�8g��f.țc���\j��0�:}�6�V��Aƞ]Q��D����;�
{�6�� q6ܹ��\à�iw�!��Ѝd�Ҹ���8��4��~��4ӽ�RJO�+$X���@1�����	�G�4��C� �P��X����4�b��>x�c�̤���y^6�ǃ:df.6?��h�6�|$�O����Pܿx���1�Yǈq��Hs�&	�䨗[�1�f�&�>���(��@y�9�ѾP�R`��Ί���%g$�G��;/�i��~Q�ڮ+<���8���,x�A�官u����PO���� �E�����́��/��ߠ�W��mY�`��΋��VU
Q�	 ��J�b����`��LFFf�V@0d�� �K8��֊��}��
���w7�y	�o���.�F��yf���'d ���E�p�6KFשYD�ڤab�,��0�/M���(�k��� �����]��^��;����D��R� �5�x��&�҅ ����Ż�8��I?>����E/�4��p�Xo}En�DȱB�݈LDMk��9�|U#���1�u9�PK�^�l0�tj���n'�07���|�`w(��{>�x.�1qy��`
��8s@�nxi�<HPD�ɠh����������E��Ia�n�y���I��P�lسSR��&�b��aW:�.bw"�1���JZ�dZf>$�$Y��	`hr���y`���gZ|�����P`G+�e~�8z�mK�'�z�Iܒ-���P�>mS��h���Y]G;:-���B,�%��+�� ~ �Yҝ@��S�ہ�H=Mb�d��(�$��+O\@��d	k�{*��D��$�3U!�λP�m��u^J��6������HcIu~c�^2��tﾈ?���FR҉mh&��) L'�4({d;�"rTy
|��?�R�C������=L�n��Y��T����� �zx�ηt�C-~�����<��z�5���6��d��׎?����G���� �˞�n��N��{�����(!%�>8�<r���."y\�H�쏰Z�/RJI9��5�h�ߦ��?����zD�k��{��<]�%4Sq9���Y��;d{���p����я>�h��oQ��i�q9kC&%\5R4x�|��,�e������Kϛ�߯DV��~�7�ܧ�/�����XB� K"� �S�=�DN���8����;�)'{n5u]<��+��٣t�Ͽ3����wa�Io���Z�
�ƻ'6����v9%���
�~V������5��ҫM���5����U&�ŤM4�U۝��y�M�Uh^�t�l 򥖀���&���*�[� o��L���O���R�//$%ٗ<���O#�\~-M������Px����N���TK jK=����-�Wr�؆����ΐ��i3!�{��|7펺i���N�\i���5�}�}�*�b1*��[	�r�{CI��W�%�,%,�*Ҭ�S������B�7�H,��@\����h +�:�oRnmA�`�/&�F�Q j  �}~M��w��Q-1�l����p�W����`�^P&y���^&r����Ԓ��$���^\�
��ƾ���o�]M����O���"��e\~���Y�^�\w�$9�y�����9(����{oe���@`� %ߣ��cW&ĴAi�9m��X1io�{����lV&��<�Hh�+򈎺"Ƚk%����o�3�����p�����V7��Z?���U� �p�8֡[�2b��ͮ���X�i�Ps��k2~�a��<��N ֣�w��L�_ш�6�qp&0�{U����A���~�mE����i�#�����!�����%�I�!#kç��mt�ٰ�-��I�1�#�ZfIt �����bگ6�L����GjQh��2�j>��$]s��P�G���P�����8S
Wm/��c��������>��o�Y�}0Ww#�KF������ Ŵ��K1@�l�a��72F\�R��'LH��<g4"���e�ǋEirʄa�����Ӗ<H�K�R��J <���c%3�������;{r}�p�5A�/�R����v%р�ڽ�x!Z,Uۨ����0󮙛�S_�d&��B����B�H���D�2�I+aL �3CA��C����<[������MJ��Ɠ(� +:ۋ�R��L�mr,H���p�n� �Ky!g��UNAݪ�e���f¤�ݎ/�>�״2�sx4dq;9�`%MT@A@��*�P�kg}��k(S�ߟJ!L�%D���3� �%1������ȹ�m�3�Jһ�N��S��%,`�υ���q�_�n�[C/c�e�c�FJ?=젥"�oˬ�B%_��Hu%�O&�k�;ւ������^���-E!�q_s7��O�.㟎�'�=ǒ�����_� ����G�����כy�V�5`y��2E6� <��h��&�R�)���C8 m�R��Ke4Yᢏq���NBbsZ�ӻ{����
�;	;E8��-��E�<q?]��2��J��UA��/��*���8��,衫�o���H�G�J?�\�af���}�lY�����A[���UB���I�r:٤������`�l_�vB���p� �-����>� «2��D��%}rO�~�%����U=Am���
��7�:vz��*��ޔ���'y\��8�����$7�jŴ�k��TjAD@B��d��S��ֵ>���������$b��ߎ�W���2K Rb�e��/�8������l�d �=�.�Sl�f>2#N�@L�1,	]������~Z��O���<�6!��.��y[wU�`$�[m_��1w�h���h3���"�T��0�h;�X�.
E����dՊ�a�O�ՍyS�ԤW�_��jC�hoPa|���o���(�=�S9P���� ,C�*�k��dj��2^-�A�����۷��l�F�q!���-�y�a/�J�;�٪[��y"ST�Zuw}TB c���w��j�&1���s�HԨ�S��:�W��j�r�: 4,u|�]?��D��@b/��o;�R(��_ׯ��7|����5���������nio�i�Y1=��f[�p\-�v��au/	�0�SL��>�+�z��tq���tw�29�|�˩�c��p�'o�Q��|�"h26#��R��1�T�����o�Au=哃�ʩ{%I�׿V����7��Է�Ќ���@7��X%{��y��D\� ��y_��aW��M���}��ݛ+�GE����c7�?���������
q��vs�0�A��F$���a��3��z�	�:n8��S��[Bj����u��ί�_[��w �烘�..X�����`h�;����8hf(\VIK!P9��Vr:11Ce��ԝ!ѕ=b���Z�#��GPs�T�I
 q)Y	��<㩫���s_���qI�3�K��ͮh�\�ĵ-�2���*"�/v���#�o�E�����O�S�g:f%rn^֭=�&/�t nl�p�  ޸"KF}��i�3TR2�]��L�&p� u��"T�P%p�4�� ���V�� d�� 8f��l��L�e��c
E����2b�I�?�/���D��?i?U˃�I>/�E�k�w Yۻ�~�C����h}|�Zt��|��O�n0�$GU�;��Z���=>?}'ۆ��� ���C�I�kZ�\궸S��Y�|U�U�b<����M�#�^ oL{waչכ!&-y6L��Ndk����:�׹���8^; �)��χ�9�Hr��3��������z¤Vl����>)��7��Aq�sa�\�L�xw����*:��/P'5�|��nߧ�~fo�@��Qɹ5[n�-5�aF������_Z<���rR��K��m��g�V�ڽU "?�(�����;6�S(F��/7ٕ�4�l�0�6>�͒헛ō���h<,�!��������MOT�mr�F�yNTÙ$_;�2PI|ک�D�g�k����
Mi������/�(���I:�P��X�W�=���4V���m��Hq2?�g�\]��%��$��#9� 5���┬Lm�p��| ��AT��zg4o�o�L	<j�~]��Hx{���w�!2�1&"Ι���䴭�nb��]:b>�O^)��x3S0p���x^�N�+%	�+����s3:�#����T�����#���;{ǔ����o3e�uо���%����4��^���#����wT;����7�����l<7Fhf;[�����A��=�9�k� ί�Ԯ2yEF��q#����I�&>rt�`a��̄���l��7"&���iE�q���y/iM�[��M�B�2��y
�VW��V�2�9a}h�Vl�wB�X�JN��s����������o�������ז�)�^[��.�7������dNbp�6A1��uW)z����r*�x)�4�\Y�^I��"a�L)���<�O$_�V��[a�-���]�.���z��������Ε�w��n�6���`�m�f	�7�'�Zʙ��!���4���'�%d����F����O�E��<����O5BZ��n!*5�,��繊 p�g�@����8���G��ę���W+��41�p���z�|~��l����M� Y	������-A�`ɟ�jjEc���^lP�V�l�">� ���me�.^����!p�R� :^�M	X�ߧ���7�Ƌ؁5&�
?����>�d���L `sl�Qox6���v���~u��=�w��a��M~��N�c���9A�6폄z�ƙr�%�>u�n������V��o�B�G��7I����m�Z���v�i.b(���ُ3��6D��˞�_��@>wٌ�!����e�<MX��� ��d��!b|����ӽ������i]Tʳ�z����4�J��Ze�R��cQ�l+��¯Xp�\�a"�h2�|�(T���q�/O��{��EΓ){��v�N��3�ym�C��_S�'c�����in�q��U������?�sO��e"�N��)T�C$�'���&9�i5)�Ե������h�\�a�s`�7�nGu7gg�k��� ��M�J;�:
=�����E����-�8uOP���~���DD���tn�~�i��;�5
�ҡ<�~����/xb�Y�m��U��Q@��v-��E�]����&�U�ٱ^}����F�L��y�񜺃=� �h7�h�+t��+���q�H�݅;�ZPHU����c�������������W2z_y�:�x��7yjex�P�u�`�>~�e#j�w�t�(x�{��!_�ׅ��T����a���G�cڷiCM��ޕ�V:V�e�8�8�$B"2��%ʆ'��B3�]��
GW4<;-?l�vlUf�}�9��bh��K��5��,�E��\.
""��b�
��!n1�$T^s���\1 �)}�'���D����ۖ�w=R�����v��MN����5)��[�����#hRH�)�F��O��(��xU�^�;������PZ@�i�5�hV���&�rs��F�O�R�F����|;�H��k�8�k-wK
6�RsJ�y��d=)���N�7��%wpk�� ���4ҏ��hM��o�u�d1P�w��O���t<�۩}ޠ�w����N4;�x��W)uDQ��zLO��6��=Y^�����q��&9l��0j ��,�-3��:��ahn[�2��:��8�`C'�eY/OsÝH��lp��p�YYHH�����}]�B��sq��I��O�Sq$��iIJ�53�T�1�Q0��	i�Ҩ�o�)���\r��q���B?���1��5�0^ETw S���FEg̉~vF~�opg��"���j1�����%$n���`�,8g||w�����߲@BB�ŜEFz��U9�Hrہ��GɄ��h�v�a��޽~�1<��U�����wQ�ɐ��0l�̺2̠K.%�N�|9���掤|�4�aH�=;g�wW�s���I�ZC�Kg,�"{�o3�!{= ����p�h3�]�8i
pD7�̒G/�d�k���<��U��̋�o\���ّ�F pi��?�	��i(~�E���w�7l�T;�顫��FŒ��\��'�ƭŕu��]�����XkO�$%��/G{��>�5qo؏W��5�w1��e�(�qil�K_�[z�YPŌ-��I�����Y6�;r�(WᱜyFC����y��m:#�����iA�`�<�)x��sk��;\;�9�K"��z80�S?�V��*��`N�|q�{��Vv
�=_���	h� �Ӂ������s�J�[��+DUr�l���_�!��&�}�!J��Ea�U�]Y�ܝy�z�B��8�9I�`����y��T>�����،w����e��neֱ-p,�8�0	,L~�j��͑��	$ύ���<1��w�+��束�dN\��)�������T��(D}�Wv�G�ukBe��V���e]v��/�t�p$�3�����x T z��JI�v{�8��پa�
�����&j�)�z�����~GE�a�8�	]��r�VR�Κ�w�%sݽ��������\�oeH&�7��^���n['7���O�f�ndu�m���9Q���x��3C�E�!��$u��{[A�����9ش�.q'Q����c��^|���a��]��������iܱ{� ���H&}
 O|T�Uc��_�䡘��@����.�����[����Qmt��;T��aS\+�I��Zm�~g8{�PTLE$E@�L+�Y_�R���S5i���������uP��U,R���_�8� q��X	�?=����r���uJ�(�:�2�If��#��Q �䡻}����w��*R��=���!UYٙ��Ƞ�i:9S?D�2O�����G�7#g������W ��G��	�����1��cַwA��ǵ��Uψ<Kw���8	��ͥ��?{ƫ�߽��m�N�O�d㭘8�;��Jt��Ib��? k)��`��U"we�TN�E������u8����$�[�5V��_7UJ��g�0結"���qg�tr���b3�O㡩��h�+Ӕ�j8 ���QẏZ�f���W@E�D}/��R(a"(�"���J���(,!%,]*
J��ҹt�"- ���R²t�7�����g�g�ν��3�tS��.[�(��V�j��G~�+Xak�F�<㙪���_Wg�&t�����4��O8�`{2�i,H�\��V_^�d��O�D�5��s oH�3;����d)[ �g��FH8��+�r�q������g9�n�����sC3��0O���)3��V%�Cv�v�a��&hE�󎎇�<����s�3�|RU��y�W��ϰК��{?|*� ����w��1Y�_ YQ_������4�\V���]�z�k�������Ťܛ
�����˗'>�)`�bL:T@���j�捸���H;�2��{W�crJ����j�9"i#�O��f�o�6�^�N��=#�;�I3d��B�+�H�ڽ�څ�q��u��0Km�r�<�x�M�Ө��b9`O��V�
�E�҂��L&�Y3��I`9PkK~�vy7qp⃩�А��`	�ڈ�ņ6���j�x !P�����e?>ݜ��}A $/nR��d)i~��b���8|o�pws���6j��t�,mӾ�������`����J�To�/�I������XѾ�R[�9��
m�R�2ml���.~���CdD �lf�83P��ų��EG��Mۛ��O��*|���O�B���{�L����l�\�~d�� �튔�d� �xjLEY!u׉�r7y�P]�j#I�45�i�*%�}�*�\�EhsH�_����䱽��
+cM�g�05��Qa�K�0�"��I�N�Z�^��5,�9e��sx &�}«z#�<d�,�zg�S��!�������sT�(�)�����:�T��w؛�5�\׾"iZ�����ZE��JnM[�@��)w��H�l���D�i::���F11�=C���l��{�6�*�`)��/�b�7�v�w3�;��8����Z����Nt�uW
���]a��y�qU;� ��PL�rM&�X�^l���s�5�-�'ؼ���g���~�ds/��rJ�X\��V�y�d!Iv��V�4F�^�0�f����q��kGu$7��D����~L�E�q+7�9�*ӹ�����t�C���� s\��0���O�5��ĵ��sqIqlF�.��zAƠt�v:=��uvz�خ�N��S�.=��3��D�7&��n�
��F�#�~l}�'i
o�B� �+H�L����.�&�5�ٌ���<ԓO_h��e2������F�u���],㪡���y"x����d�\`��/��~�u��&=�I{{!s�	irµy_Ĥ�M�0J�ub����K��E���rf����^DJJJd8%�0�M.���+����fo6�C�z�/!�ܥ�T,$�>pT���s����U��wS0�9��<Ѥ]w��n�a��ߓ���'䰌3[�ܿ~?�;s�V1��C�k�C�S�� ��$)��{6VȝF��n-~!c@��Y�Y���l�櫇�o�/��h6��橩+ �%��4�m�q	1�����|�~l?�n5Oh>�Z��x���՞D���_��[d@����ߔkkl�I~��ϢoW��4���Z&q|`�ϋVnH֖�$����yӄ��c,�û'�T���E��9��U�l�Hy>���F!��X\�C�g�@	��m�҂eI����c�jrʵ��ˮ��Aw {O6��^ql�U��^8s/��-Ȝ�+ȊQ�W
%����	*��=)�����J�B�x��y�հ&��Uӕ�c�_L>��E���^FLg���1I�i��n��G9��؇�g�dX��ԕ1�V3U�яٳ=s�b�c�`֫{�^�NF����KYʨ�ӭ6ey��i�)��=��'kG�����Qn���{����N�r�A(���s�@-ほ�+������[�솝:�d	L�BӜ�9�� ��\G��\9]�g���wn鍏����/�L�>�{�>��|4߫��j�!�,j���c��S%��M/h�}���;�6#��3�zhk�Ws��<UV�m��7�hb�"P�.��E��[��Tf�ӻ�P�<�} �*���MjfxB=���L �l���+�ȈPo�%����_:4����3H0^���c}�ڭal�_�հ��nP�ͼ���.������n�x�
?����/-a�c<���k�ks"uȫ;s�Y����:ȟ��p��Kt�u��>*p#�\�Z�p%_>)Ql����x���#ϳ%�W3��f��_�`�N�)Y{���.�(T��;m76�>�q����3`n=��m�
ڬ���|z���pc�C3�.[�d��I�HW�c�}]Yʑ5�\d(�� ���S�?28'6 ?��e�K�`=`k5�H�{v���f��M&�����ZE�balEaj*3_hX{�V�̌V(q����6n� �2Gv8#�4����W6]���lv�z ��R>N�
�b�ܗ����S��<U��ɻs���1���:ås~z�e�RfIM�cޜ��j��R�\�u�I�rr���,�!�kAP+0b�bι�������y9�R�t59ӏ2fr"(��E�W�tLؘ�쐮��WT-��lu�1U�y�<{��Tf��7���o��� ��������1�YFcƚ��C���r���w[h�X���U��n�n(��'�'�����f5f� U�q.�4{����:z��3��d�}��"�0mzpu�mO(���æDm_D\2 ���;�B� W�H���F.F����;�_\I{)���̪���˼O�]n�b����
H��:E7�˷[�X�# �
P}�N����<{�U�\�s?{y��ؒPC�<��,�&��UJ��@*%�8gv��uc�<�뗄*������a�g�j��\Qٱ��೙�����R�wF�m��40?�Cl))o�����`+6�f�6�L���cP�ic3^���Y|Λv�=��D��]���|&�Z8gc�B��F��s<����P@n
W�x.�hi���U	o3E�H��S	����SuRIA���6�=�΍�Sq����Ԫ�p�c�)���9��Q�Q.!8�]�v@_�refEj�M�3�>���*�6�l�:Ru$�r���*�!�����V��4��[\��ɐ��w�ә�N*����4�IF[���:٩�l^�F3�'�׿��	�*]��zN�ոnS��\�Cբ������:���4e��X���M%Bt����$*��n.���X�K�?��:s&��ӟ��R�K���k�e46A��zė�C#P�gu��j� a��_�����"鑒��(��þ�`��������$��_��Ԉ�7�B��X��w]W6]��e��� ;T$6�q1��l]sjC��&n�u=��צB� ���)�c�����4&��[6�g	ej܁�@ �X�ȘA!h�P|3翍hQ�n�G�xu��@��[��j2{��l9�W�?���P�L{����z�i7���Ź�H��5�
f��&؆��x
Jm��VI�+��N�����Y�����{=�}����Jٶ?�j��r,n�u9ص�#�A� ��2����t|F�T���y-�����V���{��V?+m�4NO�A?h$ L�p��U����>�m�^.�S�"�̇��LvW�Z�c�ֺ���\u�$
��6�%#K�Q dU'(~%���\����'��"��f�T�����O$kL�x�8�AUA0�v��>��u.�Zԇ�~_��D渜�X�쬼�q�]�cLeaGc�L��g�g�!�� u�e[���מ�7{d�nL-7��4�Ue�p����Z8�~�������w�� ���䜭�H���U�S�k5�T}�Vٟ����;P�Gv_�+Xa76�}�A����nD���CU-*�5Z��]"��9❁�/I�<T��>'�
���b�gYq�;��2�W�`9���&��I��C,Hثē~*�J<�JƿD�x��1��Y�{��붧�Θ�TCzu��Oo����ǘ$�j}������V�=; b�"�����kI6�V"��y��*F+������	&�� ��~��b_j�"�k����eʩ��V�ŷL.�\=(PZiHA/��?��s��nO]��R�]�R����B����)�8��;#��/�t���"}3~U��$��KcM�;�r,�Fo��5�-�ˎ:�A���A#� /d		Ji�6(�Б���N
��v��+	����^��S�5!g�VvWV2�)�Y��We`�<������:y��B[2��M����7y�����jV1v~��M^��n�^ �B�g�0�NASc
��Ӓ�M�T�ڲlj�?uڶ�z���hk>.�ڻ#�[ڨ���o�*5X�W_|�g���:u0�?_	é���v�!&"C����{�qx�A�����w'�N�FN
A�����H��#�cktwY�W0`��NBD]���0�8����顃�@�n�&����'��)=�$F�'`�Oӭ�+��ސ��i�P�� �����7�AS��m�n¯��H[������?�>4����Is�h���r�����D)���`{M�5j���N��fG�z�������\��ޅ��z��B4IA����}[�/�����K����6��U�@�f�g�
dN�\N�yߵҶx�o����΋I`��n=��r����6Y��ݱ&��<����R�{�j�
���j�����F "'bq�ރ^�(�-���H+��mS%�*�/D�����2Om�:��l�o ,aj��{�KL�[��+O9�O���'�:�Vo&ݔs2�ͣ����[���=�q �E��d��C�Z��25�k��Ƨ�{�2��� ���aH�/��� u�o�B��3�i~n�Vf+}�?�;��[�@�����ZW���#^���Pzv�>�=:z5_Vy��T�b�	qh�c�(o��.�YOX�b~4����˕��@�0w�&U��%��ά ����qj�ګ��		��q�_'d��ղ���W���p�Ũ��<7׽��>6����?�yS�+�#(��}8��7��(U7Ve�w��d�� L�L_��J������O)��6���#�[ͪ��T��V{���Mп�0��7u\g+f7
퀑��cԘgeӌΓr��F�r�e�?_:�4PE֛FΆ����K{�'���3�����m�P�ϦE�x�*�k�.a��C�Xŵ��� +�j`f�]���%�jp�)�:dc	�@��wЅ^�y������t�_G��g;�[ozj�f��U��_��G<���ϰ_��TA��59�'��� ��KJ�{���G�`��q{+��T��.vw;�ٱ
��3�0�II�HR՛>��S�V%�@�B'w���ȯYBV�g7Q��A8!P�!��q�L�K���Щ9�9m�Ӂ�5��壮��D�7���惒y�d���Զ �6�퍄E��X�J�;ee3�;뼛�S����<�P�?�Ʈ=4ͫZ԰8��N�jN[��J��Gz���o�Ō[����!
aY2�?�TD8���4]1	�����_:C�.��v�kP������K�_�Ģ����tb꣝�zFtS����H��s�җ�*+{����O�a�H��S��:���Nb����I�G��\r~�\٪j���}nW^Ch�M�jif�lɹ1a�p��i=�)^O�����'���.���W�BF� ��vk;:+�b�j׀�`P�E	a�R���Fv\ߺ$�[�|��2����N]y�Sf�rYb��C�[/7�q)������S��_�t�š���nB���lN�9��O�ĩ�~y[P��&������J���^	E������4	����ou�~/�V'����={ߝ݄�h���{��Ģsv�NǴ��$V}�%μ���J7Kw��6��a9`BRO�`��4�E�����瘖?�nOۖ�Y�ӿ��آԘ�$|���
KG��0z����5������N���c�Ϳ,�:����y8��,F-C��ԌT�5��%�������8�3g�`M=�M�G%�qu��!��T�����2uj��܋]j�6X�tb���}��x�c9_��#�FC���y~�_�U÷��te�$����pNi ��'=�m���T����J#����n����_����2�fڋ�;oPL��UmjX�ׄ�'�1җ&���w�ˋX��Іŋ��<��sخ��-�1q0f�:�E��Ǩ�Ldl����щ�1"�n�u�]v��aaU�NCI�?�9-B��S����WS@���3u+��k�L���4�b!���ի�j���S3R
��e�r�?��q �}�	������U�[X��&���BW�ܒ��� ���e��A|i��x`X��O8�Ar�D�T�#�����q4�q�w[��J�o+�x,�m�{����n�%d�Б�����Ā(��]�Z4��W���$�>��RP�K���R��G�z���i�"�Dl^���D¯�n���-5b�^�O�j��K=4�2��R���6�x�SU	C�h��̹ӋVd6�]��}�.��E8m���R&��엽 ����}���"3}�,�$�N��l�{�<�e��|�}X�PbP�/�ӛ�j৆x'��RƇ��U޷ｍ^P�Y��ɿ��uN(�!0�7N,�sF*�e6@�q�o@��÷b�<n�w�tו�Xȋ���d��������-X��R�&^�����iU��_S�p?���#��ј�)�7�%�jg�ɛPo:��e�،zD�@�*r����K����v��+�N=3�x�<� m��g��'Ei|��y1p����u�ݳg-�=K߹������h�X�����VW&�s�DGk�Vι��Ea/�l�V�U%�:��Ja��-@�OD�ϔsħo'���͡��}��gDG |�s�p<I�"�lˍ"V���1��?��G�;t�u��&�a�xao����O/�G�Wr#YP��W���$��|J�F�+�ȥ 5H�n�iE�8)ʬ�*B�I\�v)����K�<����=��jT]�t��X`r�@	d�t�*�j_ xd�DQ�cڛ�q~\3{.eTnl9���/r�p���k!7b�~��Q�#{�Y�5�G��Fߞ=��fK�� `8^p����J�}KYcO?�	��|�;�D����"=���f{�j��.����ט�����=B�P�glun(���S�|��U�YrZ_�j����KbS�o���K�A�R��.�Ɛ<��_�:#�vw��7P�$���O�}<� �7����EzMdBt�`�({u��E�%���}�&&�zV+�)kk�XƍsW#]���2['��aхnŨ���>�%<������Kǩz	��ƶ6�	��!Ju>,�_��;��O$PPup2"C�	:�0�^ ��C�].b���q1Kz�h��l��=S=����}��`�:Lx�����0��P�w8q�y�����%vz��w0��L`)`�~« ]���F@W� ��\$~=|˘�z�"qX̏���An��ű�'M��m��nm�9�y�� ���uR�ܪL��\�i���ߋ�{@��ҭσ�?.2ڣ2�	��C=in���Y��B$�q��1��6�F.�}�X���p�ϐ�~��ۧ[mvP�]�	�����aTG^�K;�c����X�B��`�`���-Ŕ�V8�*H	eC���<f6���F��@܈��wٖ�~q��G����f�4q�kw�������֎G�%O ح�d�Y%x�-�D�Q�|�P��~N����c&Ϻ�XL�����V����ɳ@���fS8�2t�~q������cs�U4��P�U�w��_j ���.C��hD����>\�\�T�Q;�z���npH|ƭ�R�^e�3 |��B�<��>��u�a�B��^ɏ�hv�G�W����n)"�QԮ/��8B-d$�����Fv/4�����J��~��LoCH;V�s����۳��$7Tq����<E�c��-���A;���hY\�)6k��C�� �8ؽ>s|�v�˓o�^�}c���*��ph��Z6c��&�-F�\����eϡC��{�ԑ�p�U@➢J -�o�"/#�)�46���}I�w�5m�,Y�1�����-���� <���v)�*���q�f�@��@z�� �J�ti;7fGȫi�U�xL�a�j*���a�Wa��5�3�5�gT����N�ԲCN~�g���t�c�a��m��]'��[�
:`�#e�
��m*/(kk�����ۑ���د_���y�bGh﹯^�k�y��<�H.�'&b���&W����H7Em�i ?���3�l:)-�Fg��	i��,ɇ!�k8
Ɏ���'�V��TSgg�t�b��]�ܯa�#�h'��z4��~�3K`~u<���"��2fa:6W�����Cl$a<��-!�z��5ם�l�[v{�4��)��������N��~C��
*0���	�g�x�%3�/+�Qf��N��G����PPU��������i�H6Q�����l��%����Y�і}�>o��S�� 91�q�4s�� ���XF���o��MVAq�kʜ@�z�܃ni�r�`�'{�@M@����4vTW{}���6FQ�Sߚ#�~�o
:����X4�e����<�=�G!�ȯ��b�e���HH���m��X�H���K�?���s M~A�����-Ó��@�t��O�0�n���W����ړm�7S��}|*%�W�g����/��G+5���̪���<�S]�7��K���`t�x�����u��|���F�.���&='߱�>�gO���!x'�`���g�/d4�:�����]�b��%�:&���#�;<	:��}ۑ��x�+"IL�����5�ǀD���^�,J;j=�nr�)��?v��Z�t��1��a�?��K�b�c��*�(�l�������v�6������{�`"b�ƌ( ��My�~�gh׼�i���%]�<��ڒ���it��_	G����_)�M5�
���JYɱ� "�շ_;1�U S�5�3�PzU��K��:��(����ͣ�(̻芩�'NiPg�s?^�I�`�MIá"���8|q��Ô�P� ��b�Ǚ��aY�"Y]�:�ٖ����a��}�y{T��S��1��L �]
�,���9Z;
m��ĺ��� T �4���֭_zD�L��(��K�D�q�G�?l��А�?���P\.T�U1E���l5�`��+�n�<�UfR�~�B'�g�9�Pci�E�/�Q�[��r���3�?���︌�����V�=�61��U�A{� h8O�?k�aZ�/�g�2�C��4k="Q���e���R�BG��Vk�x�D����}��%A���+�_��X��;��Ӽ<�ao%�i&v��T1w1��c�	�S=�:�����Q}�>����P�O���C��~.�R�t�6=�&{���^.o��z���G�@;�.d���z��xh��
�_��E@I�ɴӠN����حpm�n�*DP��'"9���Ϲ�~)���X	�	�7c/x�?.���Z9;p�Y't���i�֦��e�ũ>Q�DI7�AL�l,1vy+���U�K<e���i���6m�G�J~�ި��i̪7�>u� ��>'m�8,���k�]D�m�n׺UY���ÉӃ�޾�{9�����us��c�)�ͨт_�D�܎lʉ=��}�at~bf&��DM� L� Ŀ������s��������K����zn};�y�^��p^���D8}�ت:��� ��jⲥf�<�Y ��&�q���O�n�4�\:qɳ�����;�!��L]=n�޾O�A����]Z�®��u�����b=��4�ßSi����!�x/�`|d"��������ƌc�W�Sı䶠�����Ƴ`�9�Ӻ��i�s�S��`�+�¤z�8BGQ-����DzxX%ou��fR��G�dKeWa��������������!�I�XN����8|/p3f@#��' ��
C���n��7\L�i>�(g�M��IE58�ܭ
�:ni^^�w��E�_�}�ݛ������ȝ�h�n��2c3J��G�}�(E�e5EF��ـT�9���V3��������)X]�7Bb�u�3�⹧�$���C��� 0<����I/�~8=[vz4LE�^mpt|��z/����<�I��;���̩�wӱl���@�U�zߠ�����dP��bDM:G�H��V�2\`�٢+W7J0���R��-��.�*�����e��AFO�PP�ꌮȾ��J8���2�G_Ei�,���?ܽ{��TI�c8�+3\JZ���d�u)����Gh<i����P�G��7�ި�����ZG��>�O��C?�L�1�#�t }�r}�>�hC,/n��b��<�Y�����Q�I l�mU��ſvy��x��خ ��Vz-�/0x,���Vg�4�j|�]�r��������q�,=�#��m���i��(��.K�X���/!���l�n���~��3�p�Yo�G�����jk �IBٸGN���9��8~&�����_���y�C�ToX�,p�l%!�� ��r��C��מSi������)�=�3U����'�W����������"����Q���ܥ��D	(�n����1G��̀T����p����0��Mfx?O\�� ��K&�b��{*W��f�oD�3�܇��Z9<Y�9N�P�f{�XF���� ��W�����d/*�CْvMMA��ܽPO�������?^&^���C���m�o��T�9�N<��G����s�է���������'��z���ٷ��XF���SP���&�<��a�@œ���I&�&PQ���$-�]'#q,Q�N��A'��#�򊋽�'^��g*���n�r�K�H<'`x��j��r(�ˮ:Z����P'
A!@�~ߡ~^���s�����d��sxa��8����8�{r�Y�g�n��#w�R��+�U`�4�0���_�E���l�2g݇:r�u�_�$e��4�Ī���E��������H�Y1[ޚ�����<��y����i�/�y�(5���Y�D�Ϭ�z�1���j�P�	G��X6�o+�=��#���e�|�Ъ��R!���r���,�Tǌ�#"�?d2h�ٟ-n����1A~>u���u��z,hEAb�3�T~����T�U�Pp<o��oI`�<{�E�9�Ӫ������0U��D��c����r���n���K�B)h�tr/���Ka��G��h��xX�o[�,>�>�z0�?�����FC���T�뜪g�8yߩ��*n0�7A:��oZ:=�i�}쿉�"4n#Ԣ�r�%����bE��=�O�u'�D�? ��N�==�a�ݵvV�]T�)���
Q}h��M��֏�i�J�^sH`e鍽�]���ˁ�qeC���&0�2����.d��R#错b�t������xM��Ǌ\���b^�����_W�?[��j�sn4w�#3��;����9�1 �}8�4�.g�L�'����8���6^J����W����~ח�Dm���:k�}E��r�=i�w��ꗦ�F��:�ʞd�T	�.Z���{�u/�2���s�Xs�X�ԕ�9�����D�K5C�8����u�u�V$��ko���7�r��yv>��':̼P6M��x�x.�K�0�Ƀ�W.'�Ϋ������&��ۖc�S�6��T�ODY�ž�Cݶ�M�h��;�J*1z��P׊W�?�k[��	��}��[����|q�9��R|Э�4�r��)f<�eH��ӥ�Vƥv+��>�H��c�i/���F���ng6���`x�t0}�a��H)���ڣ�b�R���9h�B���U��}���ߛ�����+��:��m^��e��[n�(���u����ߜ���')ٺW�ڦ�E���@|l�^�J��<ڏa��O=a?K��ti���g:1ׁ��`�8�'��{�b�qy��T�^��:��ؕ7���<�3���a�&�w6�Uk�oO��n�M��������V�q�_9�$��@bd�l���~�{o4�G�]S͑՜9����C��γnQ;?�3Ψ�b0:���j=>go���J�ԩ�y ������Ȼ`�L_X�$��=/8�ỵ�'�7p]��OK����U2͑����q�`zL�ã{�[�U����� "ǉ��w����%��ը�ٰ0��H(���}�g��R�_�o�:�K�p��X�j���
�-� ?��"4�skS$P�����������?�Tθ�"��|��t(�h����首��J L�K|�}��1I9��T���!-��B�&ibb׻2t��ֺ��Ɛ�a��Ҵ�d�2&m�&J#kC>H+��]����>�N���a�B�%X]l#F/��j.}�17�C$e'��E}c Xo]�������QK]!�E�0���Q�unk*!Z��#2yK�� �ź��;ɋ�f�c��-�j%-��iZ��
�Ȣ�ǽS]-@���^�b=�@�j�?,�����`��Y#�h@��G�ygښZ���?
��In�a��+r��Eb��w�x�I9��s��8r�w!�ȰX}"�{��B��gْK�H��|x��m�F�X̊��3��:[-�d#ơ��:;m�H����3j9h؆6B�����E��צi*. ̟ս��E�8_nִ߳X[Xgbx����-I����c��czlupSi�L�����ZjsM�UR:�4��Q�_�}<��z|�M�9Xd"����U��);�=�y���uK� �;��`0�7�V��]I��� H�,g$AFL�r�ޏT�"�+΀{i�����
���.��6\'숥����sw�2r���4K�ۦ��\J �V7?��<��[��w'�
��3����H�$����g�\�?�  x����t�J-~�f���M~���b��\���Ŗ<VN䤩:�jy��&7�f���P��g6b7�m�r�b��^=�Eh�_P*Ԛ����������ح���{A�W�;k�9 ؽ�1��	�ټ��"��?+�~NG�y�.p-&`��8�� $�7��7�*�ZU�����[,)��w�F�&����D��	i�Lt���(�%����� ��ɋω\�_w+���xg�aĮ����l�1Ƙ��\+a,%tR����;B�;[zEǇ0/N�����P\N��i�P�G�y���Mm��Z��[L��i�ÙP���wZj����Ȑ@R����y%���sA(��'�\���̥�4E����U�ZW�'k���[|ν	���T��y�����Jg�����n��-�[E!n�z�zKGu�r�wLy���b4��(<����K^g�]G��)Lq������W�Kso�E�.g&rK�5T��������:�SRRAk�hG�?eT�w%�h�+L�_�����ۙ!>�嵚�z]��&Xo���讐Jc��\��`��ڵ)`�X[Th[ѹ��B�J�Z�*���T��tl��>{�Ჟ����-�H�KF)[h�;ܦ��1_X6�W/R�\��\�
%��ώK�r��L��"������vr�K��d�&�`o�������=�4g� �f�s��&<�Z��Ǎ���U8�6A5�r_�������_���.�3���cDʵ�Ō� "^N eK��f��ܔ��~���tk��������W����0�4wu=HI�л3���x������#��`C��i6��}UP׸�hV��)]_�������[��Wt�#����x���f��	}�'��b���N��/�b\�a8�G��~�w���p�U�\2f�׾�g��<����7k���c���^�2h�>�B�Q�*��ƭ��/�[�L5���?u�fi>����B�\��Ҋl���e$:87�!l�T���߰.���<�p~
�t�I��������sہ[Jr�V� x�f-6x%�p=��uxή9;���3�k��o�C��nሜ�5�2����%l�Ur����9*Fi� e gW���#��j�H3������q�w�i�O����_�w�u%BE�9���DiW ��D�)�ǧhj��a�#Y
;��%s���^�O	���V%Z�Oe�gU�=�<tn�?�������˯z4�Tn�C��ɡ��Z���1y4�o�[L�H�p��}]��4K3�p� ���r�g3�6
V��ч=2�h� �?�.Ֆ����"´�gV��"SL狼�+kk����4w&������%jo� ��pӸ���^�C`%g^"[?qT�A(HD{�|o4��e`�u˺u�{kS&le�l@� M�M��G�<$&'_͊F�	��U��~Z�
-����e-��j��tx��hi_f��H���AGN�e��Rϸ������Ts�~w$\�� ����Z`����s�tn(�#��� (F�OdQiή�3�\kt��<��̱T��M����&�ô���C�j?Q�?Z��;t_뒕�G��ࠇ`��~ �AOs�Gj4��9����	L���N����X��G�T��D��D+�u�_Hd��������.clI�3�(Z���%��.x�	��j,@&�M��,�:�Yo�;%��?hO�=Υܜ��@�)ˇ�!���.�ɵJM���b�.>�sX�L���	�����]��^ɑ�?\}���5s����s����<���m[�z�I��cW��NKxAS��N�y�f�}��⸨��Km-��5�
�{�bJ�3{��
&�'���?E"��)X�s@�D�cD�U�P������lvV���a��]���g�\S��E�`�~����P_e�x���δ��y��<+5�A��g�K�,5��^VͲ�l���]2�L@�:K~!`�����I+�~�� GI�%'H$lyk��u�E&���D�^?k��'��a�����y���ʿ�6B�#wf��G����,�zi=�AM�8,K=3}�L���=)��`?����m�'!Ht��9���m�&ȍ�ht.���g(�ʞ�(��^ټ���S5p�]��ZG�\�N�!7� >�Cf�g��<��+�ʷ�)�?8��i���p�kC�Q�)MSZ=����`��	6z�{�0�Q�y�K<@20~�������������V����t�����3gZnq��I��Al=�7#�|L;YZ:��}��n����"{�c�u,�8]!
݄�QŘ�Y=܏f�D<��!'�*o��y�]/���*���,lKd	�C sV2õʮ������L4ە+.r�����)L|=��-��M���Xh
��պ G�k:�}e��<�|Ұկ�1bA[(�9��4K��i���Ol�g�_��I	����&f`>��96�^�����9�cF������c��w�֕5!m?-Q���m�"�ZՋǿ�Dw�u�IH����^�}�՘��K?�@��e�0Xg�s��H�&���O]~�����C�t���o�&�o��!�i�|:}�"[�d�F\���Q���"}��o_i��e�Zv���x'74�W�]�~g��&$^9�ڇ�[6a�_���J���H���}c���j+ל�ZYo�V8I�e��g�}��SůFn��ߖ�"�e� ��Ng�'��T��úW� ��|�/�.&�?���5�h�g*�?E�x���P��������W��-�>��(:�����"�Zz�h���.�S���[8`�yz�L�+�4��>\��U���h}$�5��a�����+����� oNz�in�����l�4����%D/b!FWVЌ���je{M�����O�<R!_[P�^�ہ�9}�Д �E� ۿ��$��y|��9'L$���_Y�3V�����t\��޿C������z0T�Kڪ�M�����0х~k�H��#�C+��RW�FSo�w�(�WM�54q��P �'�lGD�Z -��e��FP\9�]{�������Ϡ����Vƫ����UT�6�L��q�	��&d�X��	���";��>�iw���y����p�q��Ahx� n��wɚP���Yt�m�|
�G#=�y�W!`j�;�u����C5���iD�����6g�tu�&��"d�7�\3���"��z�	� " Nɇ�P��4��R� �&E�{K�H��4(���u�t>1��*w����<E{r̻�j�Y���iq��w��E��yɮ�7{�p ���I��*5��MOG��7�a0G��?:�ݥ��F�A�
 I ?勷�V ��~m�6ȥbh����V�Д=���c@�y�i�X��������Rӥ��}��-�F!��c��ыR 4���e��u�믋0ɿ��zP6�d����}�&�ul���!��ٖU��������5�L�a:�e���+��C�psGV��j����� �*%׊'��2����t�f�[å�M��_ 
[k7�*��0�ȹb���[�](UZ�c��Z1���C��Sp��`��;�޷�0c��o�"��ϺU���ח"���:�+~�����H��`��m�9������u���⪷֤WʹŊٮ�&�0�J0����|�ù���[Y2��;���Os��#����쪴�M������I�ѽ�-�� �0�L���g�n��������b��{	�t�ţ���C�F����I�q�x6���R�j�f�	��x���>X��u{�Cթ��qj�7�VD$���2ʎ^@	���Oj�A镾Ktq���Y^"�w {4��Z�{�)�c�k3�~�����ֵ-�䩔@��+�"���_�~���a��#ڋ�T���g�xRV��.+��׹hc40_�b��G5����`9B�.�I�kׅ
Y����;����灝���U��c�|W5����v����1�D\��4m�.�R��������z�L�t�@�re$gWC���5>�����Aj����p@�P�� 5��3�m���� �Z;hob�����T�?_ �3�0��e����Y�nɳ�i�FO��L���^F`:[�Г���'�
0(��!�``fי)��=�2*!��9��v�K��/v��<1��78\�w�8�?a��:�|�?�ѱNo�>CjDA%��b�+�1������
O�ݪ1��v[`s�����f�c!%�̾��P'���}K�+��-a�bX�I�䆳����cM�|��(6�l���BP&��󕉹s�%�i��k[��J?]�v�+c�R� n�~� ��[�F֚Uo�B����>@��Kej�� ^:c�gi��	r'>�����L��A@t]�3,ƈ��eAJ>�Ek�CZl�!x������\=����W���~����q�ǹD*�YZ˄@�I#@��^w�7cߐU|�V��,jI���]O��2�^y��9�v��z�y�;�Tw}���co(��5n�OwW���lF��'P����lEV��Z����iI�>�C��ճB�{{4�Q�7��2��԰L5w�4f-q µK�,<E#��xB���wb��Ʉ��}�Oz~������f�šN"���3���0^�R�6J�a�w�тu�t�.��;��.����aR����y:�p�*�n��B��vۅ�����#uga0������ήÍz��N �ډE,|�Zp_��1�ɐh)�(�[BYW*��p�"PK&��(`I��څ�}�x�lzɨ�e����+������Y	J�ox��ЬP���<S�e�ф,��4{��t��m���Z���r��9�\P��S`��F��ߓ$��pso�;h��(���M����<\eXT]D@���C��C�N鮡CQAR:�����:���|���<23��Zk��F��.���m��öNꮨ��j��XT�j��5,���x��.���L�,Z<�eG��oQM�,�������B�_��On�1���$"ҤX�� ]���x�6����@��g�� �s����
���(u�a$���O�&�9��݁���ql6�C�����P)���n}8����qU?ȕ��`��f�㨷r���5��p�<:�ڍ�9�@�Ӧ^KY�4c�;!&�Gv�@�[�p.B�aN�Cy��-�ʥ}�Y2����c�W�(ZS&���������=�@�#�3��R~������WA@�,�,�h$F��P���J �_���8�ʡ4)ܑ�������UE��ʡt����������P�Ii��5_�;x���hc��)?��|8��F��]�~��5�K<f�� �J���F�]݄ÿºiD��V ��ih���DĜ�� +N�H��,��i,p�}N!¬������P�
-�D®���%�жj�.�54X�h9�@ ��k�փ��Xy�P�2@ުr˘=�� ^��"�T��[�tfh��ه�G��Z������]a����ԟ� e��qڕ�{�������5w�Pn%B`Y0p�;�T־6\��
��U�L�&�� �t� ЄWi�QaΓ@X]n�S�]��'o%����oM��3��s�ZI���`h3g��Y�;=����K�?t��n��U&�Ո(��xx�Uc��" ��E�\.�vZq�ȗ��#�n�%:��
l�@���`��Py��鳅�X~��ž��3r ��b«x6!&Q���
� ��g{�΄7�wt���b�H~����i+�3%�Q;��X���sz�S<E �w+�_f�py���@aK=$� ��5j��J��	���a�V�2����|�a�X��Jzu��X9�}i�V�M��v�g2�K��p�S�^�ҜN�i7��d����;y_n^�����!������!3�� ��x, -�(�G>�	?���~ǚ�78:! �\���0�8c����w��]�P���^E;�E�$�+&G`XT�^L��![1
�!���C�M h�t�;v#�~S��@ .��I`��#%�=`��i����Dɝ4�>�rΕ�.>�Gb�]��óNw�r<�4Ϝ�2�������������6-�T�����S=����	��C%��OkD�}-j�`�5г�a�̌�<-:��g��B��8ؐ���r0*�^�Ċ~�QȀ��_��v��:i��\������������99Z���t���s�4���iK����hxI�S[-K��$�
��R�����/�V#}�d��Ԟ�v�wsv�3[���Co��˺m:�S����~Q�+���[����unU.�@NP����JM��ͮ@;�J��}�����=a��&��f�3��9bv���m� ��L>/��swS�'�c7���G�f����&F�%Lu����v8�A��CYK{�I��g��F3�� 	"�u������x�� $�G�z>Z��ɰ��jA�6J �ӱ�d|�<�Z��c	�������'����2��:(}3ш4���CP��62A3���E�-��q�3��d>QXVh@�@��F�K�o��?N�M�YPpe0	`����h0�߰0:�Q�^�O>�h�&a��Q,e�.�4���O�Y�*�f�J����PRp���N����P�L�Y�$B��y5�%ܓf�i���=��?^�ץ%ǎfR�6���j�
X׈�U}��u�+>M������l�L-|o�	l�����g�I~��6	�ƺ�5˪3�������ԀH0������w�*�,�a�C/�+�w�� Q�U-��w����p��Ӡ���t�%r�n�=��uI��r��ڇ���D �h����+����A{-�~��U %��T��hB�S��!�|��"�gm�azy)4ɞ��*�f�ƽ ��r�.�0�pe+8����b��zu�z:x�b��{u��r[��jk�oe� ���_U�b^�d%����61��7b05�1N�g�������S�J�v� ����g�=*6h-!���������'�.�l?�����?���N!
iue��po�w2Y�>���a[^�hT�d&sR��lB�ȧ� ��'��Q�c�S �����#
Ni��#:�l����\�}'y�d� )\�����ݤ,t���2��1�^���)A.l��
���UR���(8������b��zqV��I)�8И�'����u�f#���p(��S]���hI��kE ��u� �=-^Xb�EQ&\ɂ�9
�� ��q���PQ����eHJ��q�>dJQ�Ӂ�+,�z�8Dt�/�d cX�Ͳ�x�5���q����?跴��zJ��m ��]�*8t�`}�JsS�W�ju�q�<��$.{~��o����w�?�G@`q~�;�{�:,�h���^�-C��b�B�< M���h��Ø��O�O'�>�zQO
�|�"#K5��1E�C��*��ů�f��q�Ѿ3a;zG���yDwБi]/�V�ڭ�\�����~?��K}���� ���E�|7�hH/�8���.����]��;뫦�`s�V4�]EA��hHzx#��&��`�����D�ܜ
,U��W:8�{�]���38�TU�d>>�y��b�$(</a��-'��(YOXl<�_}}�q���5�T|����ER�l��r㩹7��3�D���i����d"͈ՙ&�^v����g�Dw})��g e.���d��x�\0{��v�xZ� �OL�uF�H��0y�\��l�Ȃv�����V�p7T�� [���5{�t���"Y�M3�>
~����|x�^P����3�'{(����^��8�<�2EU͡�)����� �|(|���n��0М��U�{��.��+��A"
i�G�B-ஒ��8��p��7�jm���?�Ϲ�����[�ħsa��+}���
�-/�V��c�L����`qu�C~7�*0�$��.@��7f�?�O�n�����Y���:�[���X���������s�[@؇����	��C���o$���N�-V [pd<���}�[�x3��>M߻��dQ�K���0�.�b_�~�2�"����F���}gތʽ/�H��v=���l���� {� P/Uiף �����	P��ۏ��.�8��E����]Y��h+q���w��/#�����?@������������mMBy��Z�����F��K=�q4��^=� ,)� _V���?��;z�Ԥ�?QsZ�00~��
�咼��?k 2�A���$�{���~���l���[�
)�c�?��{��6��kh��K\�0� �4�����&Μ|��+�����J��J����P�#��u����L<��<P��x��(l��wi1嬜-�)i�A����v��V����h��˭�*xl=S�;Ҏ��cUmt�W��JU���[� ������!Q���v��e�iS�e��zpLl�j��¬4.>���=���hO�-t1�j���;^H-}(����k2&{���������P++r'e�F=��8*���w�6�F�N5�m�V�_�ُS�\�ϛ��r�z������$x��ċwmK��[�p��L����ݻ�]�s��C�a��iSZ}�E�O+:oz6��9�&H5{oX
p�����/��5v"x��>�e`��7SSt��(�o1�ї3�n[]�D����*���H~��ϲ��ϧ�� |U�!�%�ǡYۍ.���yn�Lw����xe~Uw�G�e'��˩�H����f��Q8^��"c&c�gyΛ���c�hgY�i���!�3Y �n��~E��$�06��0[�"����E �1���ڪ+�xO�p�%����M^qކ%�)\��w<J\�n�w���	�W��)5ԗ����K�2�B̎ ��P+ߦdV�'��}/⋻�P�)���ZJ��C����aSՖ}c�l�O�ǨZKɷ��jrfS���<~���}/���ϑ�uQ�>*��ΟH��5d����bRR�,RR8kUۘS?za��L�8�h�
N��w}z55�Ng��d/��\�@f�ШITe�P������n��Ȼ)� 9�of��X>��E�؞:Z����<*]�~s}�|7W�j��	��zV�6�> $Z��[薋~(�p�i�U���l����=}��D��;�<t�A�\�VY�Ӳ�7f���!��>�Eh��NKW{J�������gf??����FŞ\��W��ۓt��<б�
�8��>Q�V��	VE�fzE��!������$8׭o,�jX>p�X/ѲC%�J�����U�*�2I���	�]7��?�|twG �ج�z_9�ǎg2fY]��t�r��1����L��k�=�d&�u�P��\�J���y]����q����(���tw���V~�W���f�#i��Tpdd.�����om��M�����4��
��6z�J�0u\<t��O��lmK<c�߭�����(��q�P\	�g+W��"�P���X����#1��)��x2>Ńm�9�ĭH?s"��a(�LF��~���y?vf@4��un����1Y�x}*S��L�''�����!����A�
�F�V;߯��G@����b���� v��^�C�Z��nB�-&��>�H3��P)u	�����a��s�RK��t�	Rms=ˮZ"
��?���jjs���5�I�a���F���q���d�A~��� �N���giQ[������;v�S'��or���U�A8Ɍ�-�=�X���?Z(�x�%i-*���y!� y,[q6)��X"=����X���q8v�<Z݊���/��y������	%�>3���Q��+�n���%�C����w�]b�����+$j�����r�uu�
EQ+��5��F�qَԽ��1�>����E�_ib�k:魏���_�@�t�/~e(k!�{G��ä���iP�WVWI���y���G/��ٝ�v7F�T�=��UM�%AhJ͂���s�W���>!�T�L������HN
���w{��9ك��NHM��>R�9*�o>�i!m6�k��>����>���j�(��v���W�s�L�A��AM~�/����W�r3�يi���r��#�̢xS�WF ����8b-����u<͕��<P���Q�Sٺx[k���8MI���i�j��?�Uq��Gl�s0,�ʺw�GF^��J���A�hs�FSP�8@��\ǭؚ��k��&	D	��W�f�g��9*x�����f<���8��fc�N���ji1������O|�s�滹���q2���N�"����\�zJd���dD�* .5���,V@�.���?����2�\H�\����SRT'=�啕�^6�ϗ7l��!���9TV?r��&[��Gw���u�g���V�}�,L�^/=�jفv^�Щ%x��d�m���D��̭��ܾYVV�����Z M�5M?��^u�6�����~�Y�*��5d�HF#�\�>>���V��L#��4w�lIP�{��v�	���� 	��W":?�D$l���w�a2��sTO��X�f\Чz�tA���^#���-͂�Fr��s�[��%o�`4`e3����Y��J��,��z���t��02*�}���qt�{�Hg����q�o�]y�É��P����]W��ĴZ�c����nGf�<���}���H�_#bw�(M]/�yr�d��I�U��l�sx����tnH�۴m���ї�!9=y�;��s�������a��R�Ob�Aq��Y5>�y;��VnX�����6�$al����&�x�r)&�0蠥�V���SԞ]�B��ʼ���ԶU��|,��E�$��c��KV,b}1�c�$i�[�zQa�<���Ȯ���~��GI=�n�HӲ3O�K�����p����dio
��4�Lu�F����������]���9ţ.�� �P�I =�"�,��l�z�,�v���a%��43oe@$<C��-�V�3%�����%�Ʋ���֤��Ws5����;�W�y����|�u�8әܻ�ժ�E ��Nkd�j�nƖC{5���wM��`V�H+aF�п�y�vva�GKC%��ﯼ�a����T�KA�)�pF�� snC�*�6�hr��K�����9Q���(�1��,2+iH���
��͒��9u�FѠCr[����it���B
<,۪�RpJZ�W�)�n����c���K64��f!%��o�2>�`���h&f�7cG���N�w)T�{�M0,� "DENw�s��l���߮@�Ϻ�+5S��d%�I��>5L�w\3��F��]�RX�$ƭ�l���P�tLgM}$�Jz����M��"��TGB�6cpP�d�ShEq��.�����
�B��Z��gtnkc���Y-U�����n�*���o��_��U�I�x�H  ^�J7T�Si�k�۪����ZΗ��ŧ�!��9����k-�v�t*��=�!!Q����9|%���C� "����B�K���6��-��5���������bn��7�9�'?t�<Jt����\SD}�iV�48�vZ�F_��WM'ڮ���8�3��p-c�)�-��D�X���L+/t�}��['s5�qy7ݷ_�ĝ��ʌ/�JV��U܉�ۋ�E�{�|�9�`�pbb')�3sL��Ƭ����@,{������_j����(��:F���g���7
�@+���y
�`4�e
}�r���k�)�e����f($��oBf<h���ڪ�곅�\YZ+�}f-ڔ��w�C��i��N�W��W�v��Xw�q�à�XOz������1##�����,}���@����~��6��ʙ�;���.��?�MZ�7A�	�T��H������X�5�U������?������44ߨ����\UD]�г�UIB��֟[��!��y��*���]�q��nG�s�32�C��C�����ed$���K�8W�W��㎵k�^��j�ɭ��	��ThD�e��[�ݎ��^�)�����~�{;bl&7k�߉RT>��pR��(֎�z�m �;�[�+�\�4D���Q�0m4ꃏs��,�Q�R�-���}��n���g�����؄w�=���d���E�7[���?�k�_���A�4~��Ay��">��Jܰ�v��]�[i�j͚�`�C��[��|墘�bMO�ϥ"5�_,�ln��������u��RI�0��^Z��;C�y{����7��ƌ�<���!���W���VG��[I��C���/M@�AKG�_%Ռ����w�F�͔���/�tPFg��|�͓/f�>�̷Y�i�i�e
��K�-��L�(E�����y7E�s�~@���������p�P-�pyW����]�+
5i���e�Fo{7����0�LO���C���=���/N�4�j���o����@z���˳��̲���jKB��3-*e���T Ŏ��Y�:g��;�VG9DS(����$c^g��Lߦ�#�3d��%{�F����*��#"l����D�����s�g�J�Y꾧��l�ˀ�{R��Ҏ<��sC�K��(����[Y���2���O+��V(����ɻ��Z��� Y���g%6�\�y��hZ.6�y~����xGU�W˪���js�3�׼���A]�>���p�p�N���Ե^��"�;Ȁ�/��.` ./@K���,�}��=��k뢝w�����!���\ܞz�&Ü�.��ee�O(Vsg���e�7�_8��T�����Y����bl��b,70Gs��(�~�ǜ���j�+��e]��H3"��=՝av�܅iT2�ǈ���f���b�djR�/v��ǭ����v1B��U��jm���\mW����Օ� 4tv@�`��Z�i��c�j{G�΁S���pFƸ�op�z��1I/QYmҮD���Y�T�Q��c�����v��������B��;�0��jsc���(h[䜙�r��
���$����Ò����5��)�'����]s3�����
5[4�����A���Կ���:�O�H�F-�a�DV'Y��
,M��2���4��*7�Ѿ�村�{P���S?n�Mq"n;YFB$e[ꡂ��!�͑M���E�{h�̬k}�c��n?���e
�9��h�_�p5JY�
������j�U��<8�-p^�no�̹5E�T�r�<�3�>]cg�2k�*�JuY&������O{nD��Kq?b���3-	=l�7,����(e?:��;x��nL�pQ��W���o�p����,�R����5�F�8M�4܂��	��A��U��ՄJ�ѽ�n!,�I��Lm�i]	�\����������&t�e?�r���KMP�ʳ�J�ѲW�o�d�L0��yD������0z��m�����*�)�&=��,#�*�T��~uŪ;8ay/�MF�Ⳡ��#p�;��ʥ-��V~u�\�ի4ř�|c�/2�1��̫�|�UL��n����P����i-��s��Q�}����݈[#xaf�j��6��aI�'Ǭ���Z���hwp�Lnoo��W��h�֏��Ip�OP�U�m�h��i�8��īs���R��������s���d�m�c����t{�;�z�A�:�~(�/���P���|I�*�c�'}ZS��N��F�N�z#�v��ɺ�[�D���[j?���~uM�地o�w]��HIuE�幫6Pןˍ����Xz
syg��x��F�D-r�r�r[䙙�-�G�
H�z=X����;[o�ڬ���֨��6C��[��BŌ��対�_�lK���F/0��VD�R�lq�~�a���X������G�栧FL��yx��HFG�
ň[�ʇ�q��TQCx��W��┨���12��tW|.�PT��?���p|����G��8j�;	�������TiۙG_�s_�u�&Dcmw�fp�|f�c��6�'���Xo�)FEE�IEPpی����0a�u�AM���:3*�
y0�Ø�ᩣ�0>D�9�|�U�������⭟':`?��P3"�u�8E���[�����ߎ���˕_
+8i_�EUX�c�}uNk�:3D�<{6���jB�ִ�TcU���>7���4���/�
�b�Ep��qثdw��!���~DG��M�&�SnT�T���9�������I�Wr���K՗��x)�}XG�Z)�WjJ��;�n�{�z�p�`n���Fj�{�ݳ/�+����5ii$��8n��x3�}D�sDV�.��;�r�l��M��QN~kC=D-���ه�cx}���l���q\#i4s������&�1�B׋KUȂo���A�_*�����1�2��˯�߮��Ti����yR�����e�ffy泵�崴&���婗�"����v�}j��믬d{a�[.��צ`7�Eb5��d+ڷNMv�PQ{(T{��o��ռ�G$�ITR��=�b��.*���Y)�7���S�q�Gf�"#J�����ѐĲP���#<��~�/�K:��/��=��]���%s,�)�e��\�D�����m�
w!9�@��Ӿt_K���s8�q�*��#wN�)~⑗w����4l$�/7�b�S]\m��nY������y�B&��Po���,�����jP��`�����K��c�-�G	w�&�;�g�)�TCf4��=��^O�45L\�V�����Zn�#w����!	ĬFu:�"-�HSh�`��3 ����;����ZW^Ub��y�=�u��a�k���7p�����?��W�E���h��{A�����M(�r��6�^j��sOn$��n
;wJ��g�$$��|�gN��w3|� 1ЙH=0�ᩜm����'1�wNo"�V��5����ō��e���B���Wz�"�'�ѹė�Q��ѝ�ոR�s�l��ֹ��kWD�NQ߽n��-�s*p������z�y7�hw*�Atb	G�����X��Լ��R��Oj�'�v*npO�V|t5)�����Tu-}hߋ�%t:��h{��qM��G���������K,����B��\���ќ��
��Zd<�36ϗם��.�=f��+�~W2g� 鼓�9��a�t�m�J�t��Ŷ'xD<+)�n6�SBc��!BEW�)I��n���=�Q-	O��}b�(IG�m*(�VT�y�����A�vM<�:�]r��ǈT9����?Od��"��8��
k7���ɓ�Dy���5.cn�)����G;'�/�t����\62/>~��J�'��%�Ԓ����RP����)_�4��6	������ �:>��b��:Zuu�����Z~h/��mg+g��[����\%m)�+"l��8Li�*�MS�{ʞ���D�v��}�O�����	�!\^ݝ������ ����3�����}����?�+9���{d<��O��c��q��D� ��Bhs7|=.)����f�e��r96�A#���O�N��_�u�B9|��~�!�ֹ�T�3�b�g9�(��_"΋�e��8�ً}�]��w<��q�s1��-�G�g��[c��;L��XA��6�q���|w������k)��5)��Rk��X�w����`'�Ks�dv�X2����;o� }Ҧy�v�\��Z����xN��uJ���.���2e)��e;���7��T�0<��s�u�!ꈃ�HƢ�+�[w/�E���ܕ�4H�sn�)��f�qi��B��Գ��d��!�@�n�tWe"��+Gl���e�A��1�8�実O��#��`���2��U]vK���G�� �G�h`@;&{`3����Q���Lf>2~ei-Go�G�o5�fت
Xx�Y*�V�k��!���a/q����Gs�r��3,�nT���uxߛ�w�f8��!;I~�{?r�ǆ�2�����.���)�T5"�Nh[M�%�1!��`��*;6��e��_朴��S����ܟ�8xی)I	���]��G����i��-{�bMJM��/�ǔL��uT��k�;&�����V�͹��m�Y���@��HvsFÁ�iΥ>���$��8����Z/t�)a��B�������YX���ERk��40�}�-�[!�!8l'��shJtz&��m`�MiA�PmE�juJz�c#a��Xr{�D����4f�nI�˫�C�p�����N.'��5Q��>{����p����$�H��Uc���� ل�m�=�\�j���������h�iW�}dDP�^���@(��[y\>]?�>+����l �=�A416�����K 'J��A,�S}̑���ӆa��+���<W%��.y�b��CZqGٕ܏��7뺐i���K���OU�����)o�\� �����GI�r�(�ö��y����d��'�п���+�4=����O�	s4X���W.7���?�z��O���KQ�ud�����2;-�%>6oג���=E[s� p�#��
/�d��6R�'�j@��%M`�&��C�,V���g��j�K�u���n�����s��
�c���v���J�d�O�h�NT���n{�Sf�;��xd47��E�dm��[tK��}����p,�k�$���8�:vDc�z��s|xI��/�3랬2���O���o#�s�uW�L��0yp:>��'lJk&X�2�`�z�5n�Ѐ^��+�G�(J�^v��-v��@���z��]�V奷���e�4���.����nbqƯ��J%�;~��܎*6������k[V�����Ŧ_ ��y�B
�v���K���)���Y�Pyp��U(�{N��X���Z��8{�h�!j^.�9gB����x>���,!.=K0ٻe�BD��bߓr_����
Gf�x������2�(D-�Vu�PF�qi��{�#����E�x�#���,�)o�+G�������=�n?;�!�/�(U�t����a��y�Lpj���Mr����9v�НLD�ˀ<s-�� h�y}ڽ5ö���&<�/u�9}�h�rw:����7,\�h��]/|�lQ�p���c���E,��_TO�����9�G}�z@J̚5�僡C�%A�WC��Kn�����&�e�oMJş��J*r˓.ɱ3ub�d����LT��=��1>��?� 8��~�FS� ��8+P��M��G�� ���� ��|���e�q�� Ũ�[Y�}�W��k�r��C�(-LpԾM��fӨ��.0Zb�W�?�#�-�~��!@��~P*�jT����[�P��Y��X��2�:A2�Kj?�%����`�G7�՚�gߚiA�s��ZZA�w��ȿrW{�{b��.5R���x�%@��=�޽��
T�(Ʉ1B��h���#�^��o��TX!�L�j�W�1	��
��:��e���"�0�H'(����Y\KP��+�(��w�)(=-ٟ�P¥U�m���b����]�ټp������|�j����Ҍ̵�ag�z�%6��G�&-o5��Ԓu[ܾǎf�����W7,�ӕ��f�R�_����
y�'U�/��ˍ��j����oJf}A����$��&@R'���T�n���+34[EIK���J��-E��\*��o+�������배'#�������9��K_�W,ki���3�۸r�ƾo��{Nܕ�-��0آ�(K}�
R�5L���eKe�W�L=��4L_��O����fCe�������3M�6��Ws+)�_�Xyϴ�%nh�-u������D��?2�	����Q&��y�{�rs��t����&{�|�o�(�ݱ�8�m�?<9��xq�sV(h}҆?�;�2ͽ$L�33�9@��:�|�`����rĝ�S�	�ǜ�hAV���">y�@\���!�%��W?�+���	�I��N�K��r4�����#ӌkA�6p
$��R��=�`��a�$Q�����"�"���u��`���z8M	��u��W(�����{E�n�Z���N�J�ˎj�����`	9a�(ժN)�����*<4!�S���D��&���ٽ�̭�`�b)�{S{Y��N�X"!}$�-��wV}YǰD�{S�ͅQ4q�W�8*�&O$Qێ��½U7�+�dp�Y�-( ���������,��\��m)���j����w~]z;��e���w/� �,�(��md}��N�&��o��sg�� ח�2�~Y�y
s��gX��je�ϴ/��k��v.�TT�j�@�>r�B�?7�t��������:��V�I��]�1ޫE�b �͍����cMw1��m�Q��-�h�〉�,~ADɂ�ߺ��+11��Z �y*�� Of�e1����Է���N��������:� ��� ��p�����#�Co�.ԫ�=�T�6�i��	(��[k�Z&�����
�|s�, W�iU��r�Y��}�&㌹�[n��`%MI�`=�����m3�U\�lJ���|~��b��A�)�#� �n�P)���;t�F�I@7j���%�x�AZq�k�p4�%��ƿA~�֟��T7��ꏅf�w� ����/DcTlj@��f�-����
~���+۠
�{gxF8����gb�h���g�C5N��R!�
����C�C��� ��݀������?�=�2ni(8IѦ�\�[��� F�
I*����������C�?|���@Y�U�8��uHk3�_��N�Y���e�e��E�0J���{�[3�U1 ��2���Z�
��xw��_d�t�b�@7�j���7�`ʣ
ʗ`���6�XGIF�����@ɎU0aoϞ^��u�h�S�x�� �a�b`H=3�k�sG��	L���;���l�5u���غv)���� ���Ji�����W�p�&D�>l<H�V`t���d�d{�ǅ�I/�)�(t����Q�¤���ΰ�u_8��NbU��ȣ�k:[�y�Wm`@�X �����d ����쏍{43L�E�u�<����Nr"�t=���"Ey�Z3P-��=q��_�*����������M��"�U�P��O�w�f������/u�RFт-x�ڤny)�Ufb�?�c��<��f�N��w����E�ƺ�������g�v5���Q�5�Ƙ�� ��@m^,#W�8�c��&B��|��%�n8���t����O�
�]g*�Z֬��Z	��C ��*��yξ�s�`���+��C,��0'����.g� �_�f7\�'�S���t��f>7W�2���2 aS1}}+H�^x�'�]z�_t�t��Yjͩ�ۿ�v��_?#-(���3gz���E&�k������QU0n��~nK4����^����uK7Y�T���ղ�/9v3j� ɹN ��S
n��g	F]��Oc�B �Dke���X�,�W���d9�36w��e%i�M�5�C��4�Q���ųJD�()j�Quٸrsj��̛}��������Ćо�g<�e��1�)V��C��ke�R���a*�a�}o"�^F}����4Y�Je8���@?-��7|�^������F��oH������ӿvEN��'t?���jrJ ���LT���jeF�Y��Y0��?cPr�W��\v������l	�}x����J�\�������^�~o9�|��}* ��������y�^;yah����Z�_h:S�R13����ݣ{��S���>��-�	3��G��j�L����̫�s1=���}�K Ϙ=T���t䯒�"n��B�
-��e��~��s��6}*�
���d�)˽�a'm�$>�+^GD��C�N�Ձ�/�c��2�	8�B8����-霉XPA�y�-�P�=i2��]�Աǭ~���K\kt�G3^�O�
��e�|�R9�q�T���ݽɒ��r���J�Q�V�Κ&u�jrH�]��jt��O��֮���L�T>�M��4�Fv��$K%M}����!>��ƛ*�0w슬��a�)J=و����@�q�ɥ�@<�^Wz�Ϧ4�5NW�<71Ơ�RmI<��[�k���b(���@q�}|��8�&C�c^�>3R�빞jd��mN�}����# ��۾_ѭ�؜��Ƚp�$�Q�?>od��ʚMz�C����$2�`�rA_���Z����p������~my��m�쟿��'XT��^c�3%�?z�,�:�CY9@?M�CS�[7T#�@iZ��c��C��vS���v nr*m:�J
 ��=�s J�����*?��ϜME��~+4^'h��/��8��>�|@/���qS��:2��E<bg����"���Z�5���b\i���37}aw@`��R��"�,�R��y)�	��4�#���1�[jE�J1ڛ�{�-�𴯯�O�Akm����ڄ�w�/�K�g!��2ߜJ5�}����-�Z��C�ѿ�[>Pa��y��K��.��ps�«}���5����u?1�1��S��l��&w���~����{��4j:�f�I�x��ev<���;�.T*	���_
���Lߊ )�tʲ���yM(D�t�$M�<e�H��ؤ�ͷ�_�y����;D��_ �����t�_��\��}�w5(T�SO��bH�Mk�� '��8'�M�J ���U�����J5�yw7�H�!�a�Q��,�̤O�p�]�E�^��\ޯ���d�a()�^"!�^v��� ϻEn�^Ϯ�����y�4LT��9՘�;�6��/2o���һF�f`E]���K6���A2��@&r3����JaF-@�%���������H� ��z{�s�v+��%	R 1��{����g\�CSSo�C�h%!Bz�f ����E����(\߄I�<��3��P+n+����T!g��WB��2- �ͯ�>��]G�ƭ�ը�P?�`)�ǣ؋tE�["ń
`x)�_��$��ME��>S>�:�ð��Nwۂ;����{淗�#6������G��L@i����7�{�T�m��d�}�C��8YMw.���d�T���� U��
��������:�7�-l�_�ս�&S�j|��B�w�
.�*�ꨴ_��m0FE`��W��o��W3�RWj��ރ�T����'L%��ΰ"��ali�I�o��8%�h4 �L��sI��(��d�'�K�]�x��`Cm��!���V�N��4moY��d4Y��^��-�A?Há���9����>+|6m�.����H�Q+�Jm���,X����X��w�/�eZz�����)������R�ث��dS*��^�	���8F��q�R!�O����\7�}쑟�}Y6 �6�}u768'�K�bނ'Q�j4�ڙ*��Jt����g�e&�>A(��aW�޻8��"?�h��9�B́�{IZ����K(��O�o�苑��u������ͷՑ�G&BM��=�lզ�1���0_񱣸��W��W�a �Y�gh�d��i��1Qo#
�۠��������HÚ���Cx�����n�HQ^���hM5@����X��FN�W5d��tnG ς���#��$�O��7%���'����)s�b���!��f\��0]�A�-˛?ZI��bݮ�K���C���7�(a��?�|#��jO�ǫ}�p����� QD�?��o}��S�ܾʥ��UVG�y�*OL�o�X����]�IQ����H!1�T֛�iL*S6@�xbQ
TZm����V�61鿹�b\y"��&��0T⋽� G�U��^����呂�E��� SA4��ĉxxڬ�7=	�I�����j?T�藬!�`���:g�S��-��)�9L~��� H ��$t�H� ��@�H�������z�t�qF����/�my/-���*�:���S�}�=N��'*x�����ь�K6^:�}��o)<a�_8�'�z���hX'�O�q?�r���#�&=�����o�;�/�W�RU�䡛���롍
A;�L{?�\�2K���PRR�w����s�� {��!���R���7��A�S�է����hUsi��w�&__U;��C�6��%-��O}vu�9q��S�f����������� ^�5⏬���&�z��%�8��l�3�K�5~��`�	�f6�H�fW�ȟ~M�H*��mcMu?Q�V�!Y��d��5�I�tp~%��,����Y�gB�0_>��t�]����ւ:O���J���T�uTT��=>��(��4���H���Cw��)(�)����%�Cא�H������k���5.�̽�<�~���9g<�S�|P	i����!�tHw�$�M�y���1��f���[��$JN�ޙ�)H�~%8c9<�s����0Y�j=���%���ɷ��"��U�(�Y:
z5}���Kj�����jZJ� SXz%�U-VhI����3+�5.D��G�I�D��Y:Rl?)m��k���;��	w�Hk��>�����u�aD�,y��,�� `x^�^&����7C�!]��+G�bH�m�`E_;��j��ύ|}fa���wD��O!'c����Qw<3с����h����R��﫣2xE����AhJ�e���_�в��J~z�"�'o���͗�~�@�>b^jg���84�����s(Ƙ�	��T��M����#���X$.�3[��������ܖ�S�'4�މ�6l)�HQr�
�����1Be��]�ݔ�[>�ۑ�Q��Dh����6��<���RU�oy���a��85��H*}�+�@y�&�*g:#]'�n<��iw��~]<�g<>��"e����Z~���o����x��Q��TFN��-�����.�ȭ����L�ˉ ���tI|���]�!!��C{[|���&F��W�	���.�m����[fo�^���<؈\�g���|�ga@��g*�r�'/����]�sF:1;CN������
���JO*Oܠ5nd��6��劁���ɜ3�4�.���`�3��w�L�����܁�	��3�(�kG˻�ytb��s`i���V1:�v0�[�P�7��U��c�T���d�?�����^@��X���4gs�����3��RR��\�����o�+�ʢBWOy������5%RDF���Q�Y�A�V�<(�N���#����Q�0�չ	� Nr'�Z��3Yb��OM����%L♓�Usk�����f(忛��TS��M��[=�w�?3�������_�x�l}��ݒ�����H�M��_�_n^O�OI��M��D=�k�fR���K�]�h���fݦ�`�s�8�C���~��4jD,� h��7$�\��u�dg���a������t%.J�/w���9�(#W�\�F��bm�MPJ�`ة�c��'�'3�e����Kw_v�M?,��3C-���1y]�xY����~�n�J�|FL��=
vݮ�&e�/��)�C�V�g�
{"H�a��w��2͂>�MV��::�%�����&8����·�Q�z������ܐ������wl�����|��cZ��rvhk���L;�S�q�(�T̐�ꭝ��'i�\m@$s�	�7�tϟ��qd=�3�~Е������6{uٽu%א���ZA$Y�\{u6R��S�^���~�i6M�#f�y�!e���wYaL%{z�c͵`��.rj9��ir�S9J7�<p/��^��0�F��i��H�3��g�tO8����G�	q�eC������S�����r�B�,O���2BOп@E���J�^�0�j�w(�X�R�V7m=D~���S���L�i�����h�شD���j��h��1�u���P� /q-����v{��)��h��rG����Mb�E�i���8W�o�Ј���O?u'���=^���/��!�%�a�������rx$	�=����r\f~O�Q�~ck���:��\
/�}��n�-�ɼG,�R�w�Ǣ�p�\TP���c�3���Tݐ��������=y����|^�`�x�ZkĒ�;��>j�k\�;>2� N=�y���苧�!d(OK�+�����;�M�"ڸ���C����1�_���DМK�<	%����s
��a��2��߳v�{�y���xؾ��d�~0cROZ�ӴN�i
+X����Cx<�D..�J��(��7� �:���J�+��c4�+�����J봓g��v#e��t�U맏<�ᷲ���6����-�5;6W�Q���)4dgp���5�΁�Et�Y�܄�����*�hа#g���tnQj[O���]��fvY����H��#mm3<U�K<�s�ng1���cn�wk,9��C�X?���~��K�a/�W���EO]�EzojɟG��~_��h�"��@WC���,�������%Z,�9)ɂVFy���Y�[!�=�(�}?���z��tjQ��J����~��5�5�~�EN񥮰�A��Ŏb�/l^�MΗ�w�lxOJ~Gm� b�)�q�_�=�4K��1*�!e�B�K�'��i`�.�q`��y[��Q8C��،�'�V�}
*�|Պ�[}�������S��К&#I��%����*�K�6��o�E+fn8���s|�F��r@,�d�}���_p��F�fH�,��q����k9�C�HwX�O��4�tC����7���W.�q~
9�e��gzi������	kT�7!�U�N>�ǟ-��AfzQ/u�^��6_`�_���dZ�� ��_CrCADwy��<��<kcdl��V��U��/~Z���o���$*r֋�������Z�Bd�o�o�-l��	���w/���s{f:Ѿ��´>��B�����2��K~���@ �ȵP"J��Ժ�-ϩR��!kv݆�H�l�T���n$ö��)������&T!���X�V���k�#:![�qO� 1�@.���c��T��KJ.���1�l�`�wW���k_�bاݰ�zW5$ˢj\�qm�m�����<�ܔ�w���WR� 	���iN��7l�2�k3�Y�S"�[���_�@���k�B3�S{K�r�`k�@�0M�/jkS>�Ǖ���azY1l�7Y俩˫]��m���1=}��� ��m�P�+*
옰d���I�޴���m��u�`R�K��.u2p��jW@Q~��wz�]�u3�e��jc@\Y��6��<+]q�<N�U�Y�H�m�~��J�����5�E�����8�-f(�;�%�I��(R=6�4[>��q*�'#�o/�﫡�J��g7��(^�΁�l�+kX�N�^��T�K��ի��u�R�IA�qE.P:i���3QG�q8���)�6�M��<�E+�Z�5$�X]�--7�Zر�������[3tB��ǋ^��#b K�{c�e�{�u0)�'��v������-����5�������6e�����K֎��켹ї{0?)]Hk�����uZ?����Ɯ[?�sh��z7��Y�vYܐ�N�.�ʂ5���}�n���2 -9�t��zր̅J���9!tdE`}�]e	E�˃��"�VL7��Zm�HzZN�f�WWH=�����~������l��Z�`�����#En뮤���/_K��t�0X��ƕ��`�pM�!�J�:ԩOf�F֠�8&�nD�V��#K޹�Ρ7�����m"�Zb5��EhnC�J	[O�e�:E�M{�2�?#����}c��:�	z+� G�����U�?���@I�s6���>;3�W=�u���$d8����L�c\�i��[���M��hw��ܣ�s����'�>Hp�����y�O
��+[���d���q�7�A���:fP�/�{􀮯�|,��%k��f8��d����.��8!���ۘA���,D��q��f(�� z4Gր-T���V�� DY�lB}9�por��Qt!@^�g�b6��f ~��&֜��P�5E�_�Vh(@��/���X��W�iv�n/�a�q���%9H�����,���~������˳�ź�YJ�8M0�g��ǀ��iE�&�f����f�OJ���A�����ĵ�>�z�J�c�Y3��*S@l{�>�g��K�s-�)���T_[WI���k�b��w5��:�vG+P57�:�6�ŔZ����Nkⴼ2"$�ER,7v�+�5�"�I��8����N���!u��yEk��WO������?��}oO�|;�<)�w����9��� �������n%.���)aI��~�D�$�#�Ks�����$��ë~F���5���#>�>n�h�)9@ҙ�ȓ[�feH*�ZN0� >��
A�4œ2^���o��N.��Gj�a�b]�@�5��iύk[�̆��r���ٯI��i�CT�hw<�T{B�P�Qq�����FHԺ�Ȃے3�wR\ .�ص��a�J���Xi��緥`��;���8��j�ђ��I?l	�]��w~�����<�ne�&�� �!�g�!r��
���U[�r�[.�5�X�\� ��:QD�C}-oNd.���A��9��%|8q�h���H���c���8e�B�Gd��<w��4ˀ+���ۊX�>鱥�~�W���QZ��b�
��4�O�ͯ+WI���a�.�ٍW.R�悻l딫#Cy�]�{ö1"d�xD ��c�LMAn��R���#
?��*8L��QC=��峇*&�pq*�y��U���&f�Ja2�{9g�}:w�Ѥ2���}���k�� >�c��2�?/��;�P�[��|^L	�hX�~��n�
�����'���t���i���ؠ��%o�s∽G�m6�*Y >�_ym��a7+�E��!	]��婾m�:�.K����
_S߲��'}}\��NR?�{�.v@M]����U��_n��D?b{�����YZm�U��2|�A�`Y�к&�dӞ��S�%W�oW!��ׁ�Hl�\��Ť e��CuV��R����s��q�]��A�8f��M�$��[��J���ot֌�+-oʹ�X��.}�^�x}ڍ��ߙQ���sM(�9W����y���S��:�w�N�DG��x��]ih@O?h�����#���5��G J�t�i{���~�v$i�\x���}�~C��
`K�16��g/�#�;!����ߓ����~������K�f��{B|�qh�k�/��
�3οκ ��2r� ]�+�0D�������S83����C�~n�?p�)��M<ǟ��u�A�¦��ـ	9���fm�f��+��`�%��Ȏ�o�}����D�^�#b?|�J~�DK�������ʆ�s��*�8���p�;�Y���zKg� ��w�������!`��!���t����0��b�oi���	Yڜ^��&�*�Π ��]z�؇u*�bf�����-�!��Ƚz�RP_�#�vG��Hw�������ŗKd�֬#j���'l�d�z�hH�g���|%�.&î�������zU�/d�t��F6=�+2�v	�⽪�JQ���[�vP��q�_����_�[~"��>oSRf�T��]��\��p�$'_	�HYJ�W\Qq��^����m�r:횚j�À���&vJ~<\~���pm�J`y�RSvODV�-���:oI���(�a�7�Zk�"7X�}�~��Ś�~�8��m���/��y��E]ӗc��C6�����M0��ع�Q��{��V1E_2�\�x�&�L�޻����grzz�Hâ�^�c��L��MN�%�p�@4^�*������D�{AT]%l�M#I�U�/^/O�óY�� i0�s��9�b�: H����2<�����F�j���H����і�"��͛�y��_��\� ���ϡ��\��e���5qh8�B���Y�	/�RxA�E]�/պ���W�E�L\D�V�T<6��GH�>��öXd����S͍�~��|��W����yK�^(T���L٥}];��g�6x�g��W���p���x�|��#�C@6�J�g�uS8z�=��m��}����,�G���$�<����{��J����$�_��)]/m��p	�.��z^�٦Z�PK������,��h�U�T~ɐg>!3����`��o��U&aK�v�\Z�,l岼5�^���*O�Aqq)i�߆l)�nV�"��x�kK*�YX�tã��F���������l�.����d��������^��~|����4��@��)2Q�����T3K��H�<�z�h����ߒ����KTr[qﾝ�]w���!?�-& /���ۿx^xn��S�a���p "՛��H�p�P�XDvZ[��d��[��*�]*������^�����7��8��#�B6}x��e_u��l�>K��?��-��g3�%P�o�]�7o�n�qgt��Ҡr*�[	UH"#K9�wLWx�ȼS����RΏ}��\w��:QͯE�����K{���$M��ȣ�Ջ������gU�(r�Z��lf���j=ʚ�2�s��#��ق�F�W�~.v�ڑ8�?L?����.8�:0D#�.��Q��$NY��O8���"7�'d�*��HVY?Uʒ�4k)7�9�Q���p�}�2�M/ ٷ��N��R�}l���!X����}�gp���aỸ�_���)WW��z/��ڀ"NH�<�C�7lFn5|�\ɍmmGq��8��N��%��i�U}V�L���|���sW��6�����݃t�~o�P�o����/�`~�-c��:I��$8��y"B��5��M�8����	�y9Ҷ�l[��ÃR|���z��4�񹽐��1oaB_إ�P��\�I�\O!�2"�w���Nr��-��,۟_�6ŻX��C��.��/����B��KK/��}v.�3��8���H��FҠ󍰾?f���}m�ێp�4��/�:P��w�F.�!;����P@��";���r1����˝�blt���f��a�3��3!ELŌ�(� @�~�&��렿q���&�q�9�i�ܴ��V�-���LnO^[�"b#���a�ڣ�	�� ��^{�A�_�PJ����g��R��B��M�֞Y[� �W��q6��+
�+�0�����P����������M ���֯W6��p����<*�^�dT	�A�H�F��PY����G��^�=⣜{�d���AV�Q�c~��u����b`��C��B��J4�"#�C�h��$���_��uV%���^�!v�'�?ЈpD�]Sԓ��jj��Y�!+�[���c�����طSY��0���6��5
��v[)���x���?�;MM��w���V����$I�Wd�O�?��8�!�����uk
N ��H���G�Y��-�xdwP$-��2�|l�����o�¥?�x
��\�HAEֹ&�vw��:_+�Dd����e��v~��P�o"�����é&_�B���~��N'LO*�֠$����8����_�]*�4�������YE�%O�f���7�jB�n2)^�Ԣ�!�?��z��Mt���j�cO#���D�Ǆ��}�}�����3�9��()�|i�}|������݆�N�fL����X/7�������??m9t����Mm��1~���9�򸲜Ԃ/f��-�jTz7J��{,X�[|�xQx�&��߽̓u[�{�_�S��z��}�p�����p6IW\��#6���߻��p�������г�F��wx*�/W������nY�����ag��/��z�WH����Bz���r�t��KY���pM�|���r�!��v�\��;���`�qn�K�yP�>�{:����3=�"L����M*����_c.�u����WK>z���K����zӗ<J�Ǒ.!m�S�����f���]���K��%�4ץ���w�U��ly�)��k��C��n��8��c)s{�=C���!G罭/BQ���w�����d��k�w,+d��N��h{u��v���	�V��Eӎ��f2�?���R&��3�B=���BV��ǧ0������Cu���v�3�ip5z�n�Q�$���C]0��X���̍����nđ��9�'�Ւ�e���7I�H�`,�=`�Z��?}N��V��3�9��um�
�"K�*Me!�q�잆�m'͇"���s�Ƹ�:\2]���x^�0��aw7A���:ڟӟ�rYq��K��CU���L��5\)�s��\h^���I��J����Q\a^����`��y3�+8NL`3k��hX=Y"�T>\|�	]�mG�:�ͩlE��4�1/AF���0v�ѝZ#ڠ�z*k��[�`Ζ���RZ�{�:Z9��;�%��!����L�RU�D���g󝉫g�S����P��զ[��Ǧ��6`�6�;�֔�԰��-V��g�4(
�*�5�c�T:z�y&�����O��ҭY6#k�GzZU�{��� �@g�cs܎�KJs�P�����U0n~�^$��#Y��:E��;�����*g�x�%G�S񐉆��)�5Ƈک��%�[f��o�e��-��VW�[x
�3�'_vY��T<���,�F��2_�R'o��$Sl`����s��r�`/�O��7:8),°���#��׆�{�"^~P����*j�Q�ꩦ�I�+!���P�wW���t%��Ab�j�!����#R7�͆T�z>>P�����I����\^V
�Z���;�R[�!֩W�w񇳝�����+��g2�b�};�7�"�&��
%��u^Ql/�����LՅ��~��1Trs�����E|OK]�	�1z8gZ�ʔj���K�E#���wc�/�k
S�Z*�|_�{�����Z�{Θ7 "�/��e�9吕���ul^\HK�C��&h+�W�+�o�Jr��\O3jĸI��{h�Y���'��l��P4\K���\�>G�a�[5���=��/����-΅�9k�io�E#��j7��w�_O���̽%���u�!��( Ѝ��p�[�׆~�@z��;�6EC�2r�?>UԜ� RV�6�?����Y�tO�E�-X����̱s��ϪX�b�@
�J��f��P�G���99&�l +�IYd�+�zZ�_�y���/�$o�t~kB>�R?��d&SKQQ��X��E�U�� ��ѥ1��5xٹ�p:�s��|���Bx�)y�L�����sQ�sp)ǻwb�R�3da���R�0�i�:O�s��4�Z)�Dr�����D�B[�/l
���杧�����P@>�J_�3�M�JJ� %60�/a���|���s�n) n:�+~�u�G ����O���k�⴯�p�((�l����6��?F�����B��g*�=�Akdr�^ ���^��|Xp�V�K~;.ּ�P"9`�s@==��~�D���u2�Ձ�3��P-����c�+����{yY������f�c9[�C,m['�ˌoۗ5z�/�����p0�<D=�j�*�է�μG�!ok��t��Y�l:jd�M��E��P=��`^r�E��8�C��0��z��Aϓ��5/ޟ���'�������| ��Y���#�Y���W#l'+Q����zy����n��i��.���8��Tr�Q�E�^+�
�@/���nWrug�T�W�Jl��c�Z��a���b8ln%�p��^DO��y�t͓�Om����\��Z'6ئ��o�<����8���\���x+Lݷ"���0����8��7����:�]�"�C��s�t���j'�1��R�5ڌ��EV,�4������0�]���]3q*S³�w���~��n�����Ğq��C�ݻ��>{���}��Bfs��}��Dd8�:�B�r�ڒ	���	F��]y�p	��z�i��8�����;x!�I��0�i�R�iQq����M���1���h���qI�A�4(�)�$���2& A��q;�|��9�a��9N��\�53W�/W��u��O��/~q$E�d�/M4;.����?�ˈ�� �=���ѿ��P��%�&�����f�4�18���)8���𓛸��MhI���q�w�Zlf��:^G�j�k�[�R�������+��ݝޓ%5�A��S	���y;n�;Y�r�E�9�!'�g}Ь,
q#���Z��w�����Ku�(겎$��٘��i{Dj�s&�'�k���?�w��:drA*5,� �nj:6_����@�B��N�y���S\��jT�������b.��2��c�q׶qv]!h����"uѤ]۹���Z5Zy���z%��_�����y�����9�6����#�1d<m��f*��� 'u{ �Xim��:�WC�h���d���P%Z��W��Ω�+}���YdE�E��l����V*�ߵ!�O����ӥ�K>���I���M#��hrs}�{��y.����W�M��O3=U$Dy}r٤�b���K��r�ёf2���c�G�\jэv�b�Β��"Ɉy(���+_R�]��1�H"�J�ڙ"v�|!�Dv�Q)e�?��y���IS'J�ܣc�j	�4N�Ms��;z�-q�8mA�࢖�͊��iÇ�L��7�W�ٞp�r̕�{ԛdP���Sa�̕'�pb��������]��s��=-P7���x	3�RLޓ�~���8���V��7L$�{�5Ar5A2���m�m�Faɀ0�*��ń2��	�K�'��3W���|�iqQ �&AgAA������d��.��X�R��4Z>&�|H�E�]�4ᙫ�tV@��^8.�NWq;�"^�����u�TI�k9`�n��!�g.�w�����I+X:V!0�-,H��Qq���S���+s�V�Ã�P��Z����wS�[�HX^a�
�_��ʝW���UY(��{6Y�����Ib|wf?����t���ތ��&���V��~	�����1�q�C|�0�"jC��UZ� 	K�)��ջ8���_����5�W���\��xi��ӺMB�G���v���	Έ��p��B,ȕ��@���N6f������}�h�k����Ǩ�ȢDΰ�b�`��[g������l��e�R�M��#���x������X���U��v{(�ڤ��=+W�u&\�w���QBh��d���CY�Fo�ͦ]<��=��N���,�q�;STa���y�s������J�I�4Y2OG%����/l,^�Z�^���2¿�1���«��h��6����>��l�l�gk^?�Xi��]�4�Jߛ��5�9?o� ���H���װ|�����jN꛵s�S$'!�[C�0D?��M�&3�J�(��8>��u���z.9���4G�d<�%CN���sXA�QPTV�g!
Gn���1�ż��r�C�����=�\��:瓺:iP���O������g���_��3�ӿ�zv�s}�VR�v�"�Q;Onj�T�Q1X ���� !�sxA�Md:nF����Ռ�R�Z)��}ﶴ���
��\��a�,EO>ਇ�*W&�{sz�B?���R��6c3���I�z�bu7Y�������t���Uq�Q��Ϫ�������YK����"�|2VA��� ڊ�6l���+�-v��o���0���A��}�A���ڕ�o\#=R���7��I�R� o�.h��2�<����$=�u�\���6����?��yoT���h\&_v�E�a3}�X���}55���T��u�Itˬ6I��}�h�~�3�%S����f�;j�����ٕ�qi��;��fm��_e��^��7�&��[�w�Hί5���}�����̕z�,Y��ci����8�Xÿ��莖p4�L{Vn�v������s�%pnB!:T(����f�np�FR��<�G���kX6�((g�'�����:���� ��ԁ WS�[[���h��a�;P�����_�вZ�B"oB��F�5��c���װ�c�݇l͈�X7>����8�ȁ�R�q�C������f�[��k���ˆ�8Q�z��rh;�eB��	�a:ڳ�F;7�.���>g����ןo�^C�l���v�`ZT�,	^��qǌ[bV��C�;١9�qlU����k\�$�ԇe����Ҕ��ԧW�
յ<���ff��<t��7�����C5����PS��wz�!*ULOg��,`p��޻��n����3�t��q~�y����׈����lYR�]\u���k� �VL��j� N��` �a���f.1�[�{C}#�����v���ʧ�a�@���k"Uo��A�8���ݜ��)��a���x%�	�IJ+�Y��Cx��z8�	�Qa�N ��¥�Vj�[O�e�-��8�6I�f	ѥ��g~��W�	X1���|$3�w�U�Ң1�#6�1j�1�q$=WRd$��0!9����V|��6? +�M�3�~z���ܥ6�>�5V����vW՛��C�)"�%bv��LPQ��[��J֤m�m�J���Ŋ��&�B}��UUV,E���]�s���0罾�����6Fb����+|Py}AT4p�9���'�����jP����+R�ˢ�?w������FK��lA&�dB���ɕ� �U���`����A��Ӈ�	�[K�����';f�-���Ũ���zf�h�Z�ߒ=�a4���uu�螯���D�cM�{��X����,��K���	�DƞPY_<q�ZP��]H�hߍ���%r44^�-����r�����Wvl�1Q2�5�O���K�X��}�|��E�
�]9�*~�;�/m$A�ܯ�s��|ٴ��Z�iP�Ϙ:�_�n�^e���j�����ݾ	�n�9]�MZs�y/�P��B[��l�0��`G���ӊS�W�-˒�
ş�Y@.6I'��A�FO�څ��^���T� �`�}I.]z�/(�����^Y���p�y"��u��P��~+�c%è
y�`� }�5tBs�L�#]@IӰ�����Q�&,�#�_2:nL����<ޅ�U�N��Y�~��!ω��@���c��4��.e~����`�]������������*���X4��K��on8�7<���6��'X����ԯ��߱�b?�6H�=�+�e#��btZN2��:�o[�����c�e4���f��9������zK�s�D/N�&dń�Kl=N
D�θ�7y]����.K�1k��r��b��^��i93��Xu��c��%b�0��M���ulr���!��|� QPXV|�j"Ӎ��`��^�4�)Y��L��O������\K��g�a,N �_�=�Ҷ����:�='v��VՃ���`�e|����&$d�质g�F�kf�<���8b^h����I.wJoѸ�D`~��[���������R�=N��uehi���9CR�0��I�2�w�^�X3�Y�m�	�/�\f�(����,�)/u��=���E�!�]�|��ޤ�_�Z�]�V3Z����Ia�a����^��g*�g\m'תP)yqO.���Z[k=�����S��ʅ���J���}��.��]�'�����z�ᬜ����G%���D���o����Sd3����2�"�9J�/e|��s���B2�z9���.p��X�E��ak� ϯ,Ȣ�������,����Bo�R��o8>��6�^��^��\�A�
3�}}�rYru)��<�Ru���s�i#A�~S�W�I��!b��������Z��+���� P����;w9��b�>F�Ŝ&i^�����W��e^���4�?�m-�-��[�r0k�ab�ޢ
�������G�'X��d�� et~��H��+2���i��D�ؐ��>3g�H>�G �۝ȓH����򍚻�D��ovR{���dֲ�bbB+���ԑ��24�À���7�,?W�7�+�,@�O���2v؟���ǎ�i��.������j7:|zH��H?�ܻc�=�2^�7X�K�;�qL��ʭ�z�G�ʧ��[��Wg1J��  ��-0��uI_������h�b�4�m� �ђ�cu�qi��ca��������j�S�O_p71�r/�1�x��m�"��7=G��,؎UK���]>C�y�~Ó���_N�w���2Om1@ A�v��gn�怄�>�h0��4ZB�%eK� i`'|Z�E��qL�[� � ���^9>�m�[�G���y�`��k��Ak��)���*YO_ �fw��)/{�y	�H��Mt<s��&�?�4~��.p��挅nL��̾�����1]R+ ��^ �n@y����Y���'v�=_��@kx�|R�Au���L�nqt����p��E����ppS �?|��,��}���
��XM���QT����_qB��1��:��5u>�ۀ��?�B�t�#;��
tM95@��'U�V�i:=�ٲ����6K�t�E��Fh�N��6K��ȳz�6���x7k'q�������D�K/��h �F�%�#_K�M�3R�0m��$�0�'���ɂ��2�E����@!F�8W���<u�w��lK#��	��[큇@��� vW 벒:��n����c�)A��g�O3��[���́�@68y�=�53�(��( R��B��m��dq]�on����z�p����C)9�Y��l��Z{`�f�{�[X�Fj��@��;D\�*vЁ�RH�����O؎� ��΋������}`V�FR	J�P@ ��Q���Y+z����c�h�# ΍�q	��i�\D�	zz��	�`�bH
�y��~إm��!�FA�#�\X�~�D!��,�T�tf�{C�@���������Q 2�p����q]5"һ1]jl���W%�x#��G�bRvì�U|�q<ewv;3�O�=�� ����.�VL�a��M�b��jl�X��Ѐ�l��9�`>�r�R�Ka�fh���1r*T=s^��"���I� �:퇨���T/Yp�s$3���\H]��N��J��s����v����J��>�>F�c��2�z��?�ktúK>6��tO��Gpw����c�zΐ�>6�|���@�奚�Ά�������+�w�D5?�s�\�� �p,]�IF	�Ë9��UxR-����{ CJ���,�[FO�Ѐ�}���I �4\��l��8�w�"�$nX���;�	4d,�V�z7^��M+M#d�zn��I�Pr��t}����BP� ��(˜�F� �x��d�+����t������כ"��<�f"�5]/'s �5E�D�������ɑ0��=�5?Y^����" (��|��|�LC�0 ���r�G_z�*��"��"���Td���F���].-����~w�W�! ���C�jFZ<�FJ������M�ο�&���P��N@zJ�^�Nz��Ao���6!ۼ^����!)��m�fd{����4��?�j��}�HWEG�?
�I�5��ij �~� >u���Ew��^6��uq�B���`�e��"��7s���>�x� .�ר�� )R����B��$��>"Ý� 0��Cl�E�_�������j��9�C%E��Ay0ɛ>ϫa�f�4R�*m5n�E)�o8�dV�1��i�ŷL~u>�0AQo�Sp�5�����&����?Uz]�������z:�E���os�)�q�/ ����b���s0S���ķ!o�ؒ���`:ɇ�ڲ�@x�E�~vW��Ğ5���u�-Iy����xa��Z	u�Q�����2;U�ƕ�����g���U��YK�k����+��RϬ��'�?[�l��"�>��N<�'��J}3�8��"#��N��!k�+��_���Ɓ�5=;�7q.��Gu�Y�N?�<� >�S����/4�;�cu4�\yY�C�� sK��+i\�BF���W͡���%�=�#��K�4ӡ
����`*���$�3 �_2��Je���C
M�s蛐l�g�ygV
�����O6$�ӑ���&�3DWxN��:a*���!�`>�b�!��A�@���&���饏�?w��0t&o���"� �3�|��%�~G9D�P�d��;�9�� ���k��U���	�`������ޛMG��y��F ��j�t!e�t||ɳ��@a U�Ò��!��/�l} IWے�3*w�Cj��ϫ���'�9Z���� ]}�nMm�/Q��9�5:�n&�LESAr�4�����mFރ&�N�V���P���|��=���}�']��W$
���]��%��"��cb��J�Wc���)�����GVKv�I:��Q�<�C�O�������p�l����0+�3�[��9�35�M�!W��M���-v$�d,���@?�"���$/��A�I�� ���@���0��Ϲ������y�A�N�������J��$`nѪvs��g��=)E����|R�B�񚷄ֵ��:�'�Y�C噸�-d7�|�� ����.��5�(/�+��I��}�?���|'p1�Z�l�n��q�<�����������z����6ʹ)%�.���j�+��5�&6q*�C����=[��))vP۝�Ԕ٢�n�}$<�ʘخ�"���~��ν��۽Iw� 	P�K��{]x�H��*��2$	���#	���l95/�L���Q���݂�`��^��D���@ <��[�v�qWGj��*IK���@����\���� ���h���nYЎxx���(L�xĳX�k"�
�ÏHYb�~�d|��ë�F�5�	�!��Bˠ�S`}+ W�������$��R�b� Ȁ!G�N�k5R�wZWZ�g_X����ٺ��_L��V�;!�/A�f&��_.���xjٛH̀<��ǃІ�b�^���8��S�q�����O�
�!7q^��S��~}|���ϒ����v�_^^��w��@N����'������>��+?�I��j7��/NV@꫻fѕ7ϒ��R/o�z�{ZV� �h} ���\���Yc8�d\{jTN+Kmӻ$���"�=uc|�\ 5�ӻ-�xg����ߞ@�m�*=���$�\vv%5�� I�O��	g ���y�8��"�??m�d��7R�� �wmj�C�ȿ*Ŗ�Q=yc;��@�a�KwqL���
�e=�Ժ��C��j�;z[�X�$�%!B}�S��-  �.0z�a�.f =��^��-�4�B���Y��_�j����v&Xaxg�{�k��mz�.����߼�Sz��4�5^�e�N��|
����[��%/���������*{�w���k�
�J�()��+!5H7(�t��*J0��%H��H݃�������/�%��<����9�:v�
�E>��`��:�|p��񫺋�'��k|jK�=A�tx0�Y���~b��^*jZ�CSS�G�6�/֊ 5A"�CM��Mc&U�<tϗk4�Rs��z|�d�^,�G�?
��zَ��G,�q��8�6칥)�6V.�[%�F�\����[�@X��*�իk(��k��R�}p� 9aTH��о��R�x���b���ܱ
�0�ڗ�Ap�q�7/�fN=ɍ2��3�<�
:Cb_(�]H@�{%�J8k���$� ��B��+�����\��ҵ����|Ќ̚����a	���/g��٬/L����K���M^�Ҵ�E㬢����!hy��V��������rїpr,7O���rj*�� ���7�Mg��8�4fK�4�׌�/����]Ys��$[[ȹ��+w����\.	*g����Y�ad��	k���B������A��~����.�F�K�U"���6J�ɥ�h���,��+[ˏ� w�D���k�y����0���Y��9�� 4o�
�Hb�z�<�PZe[S��F�4�%��k3�i=���l�`#�h 2ܵ&U�3=�����Yz��4�Ȏ���X��E"%TDn�yN�l��-���d�"G{0��W��'������4��@8�ö�"/��i�FJ�h�x���=rTp�h�Z�Z)�)i������}0� RW4�L��?J)���4��U�����(�B�)Z�Z�`$^7�i�	R������4w�~�"s:\���-���[��g��Y���K�{J�����1���7��]�ӊ;ߓ\s�tp$!o�ǵ΍1n�*�mEB��#�^�ڐ2*�q9�[PA��a�U-�-Jq�k}��,�cڻI�p��a��A�ݥ�7�k�2.��܀��z���t�e�x�h�u���J�,(X@�?#:�o=�\{�*�.��ʲ�D����T�`����̷����)���w?��kqK<u�dF�0M�<O��pd��S��چ^���A?����s���է]m��{��&,j���>�Hnj�(J>\-�|g�tt	�w��:���U�0������"���B_���n{��<5����'�ٵ$��yy��F�+��}u�����6��3���@��`rz,_��yf��P=0`X]��kj��Z��V���O�k�#P�j�e+9�.b�Ƞ����L���Z���9��|�tS���(��4cLO��9��?�*�mE-�ѹ���B�j|���`��a�1y��ޱ9���^�sVj;ƺ��|P�Z�,/�т['�?�P�V)�L�U��I�Z7�jsX	k� ^�{]\���	/���p�#X��>[�������6]"��`�������g�T����{���G���kn���3�ס3[�����继>���ꖥ3�1&zYS�J���&�OL�s�-*��0�S��Tp����`��#���o�j�Y:��x-2�����w��#"�����nj��b�uf�������9�J�w�.��x�Wzf����&��Zu���竤w.�a^�i����ବ�N�xs.��9��E��k�Zڙ4�l ���>�"
�xz
>@�Z��Øp�,���l◡����^ʠ�,\�e�uǶ�Mw� im�$��?@�_@,�w7RF|(��	��I�����|O�0:y8ͱ2��ri=2lg�6��s�����!�k;� gQ��T|�v��We��h�[�j�C��k����*�����D�D��ރ�*�q��
�UN�nh����
JP��̾{}�����"�j��s����-�vZ,-���Qj��_g�=ƞ���(�=��{#:��*�O�4��I�:P&v͡���\�	!~�7M�%V�R�V�!����_lL�nӲ[���S�~2ʲ���+�����#l?V��Y��{\4s�Zr���$S2��H����ܹ���r��>�����ˏ5��F��r�����i:*��bCu�-�L$��:��,���{�}Ò�����H�������Xz0�C1*�3��|(~w�����T��d;�'$|��6|�w��6�#Ԋ|hC��AW<k�hxt�exjnlڴ=M�]7j�
K���.?�ئ�:������v����pc.sG,��ˎ���>��Y��)q�`#S{�ڳ"V����/y0�j��f�?aZ�Щ�S�c 9��X����gǦUhGd�yi6�
��]��{_��f�zT�����0��m�{y�o	ݧ�%ʡe�zD�j��r���m�l�����|}�_x�gN&�C������RV��J������I����R�<j�{�J�R�s����U��Z~�QJ�����+槗!�����V-b�JqRt�C���Y��I������8���<q���B�䨶>.�|oR��Y��8��Ak��H�m&�qK=fم�3��B[}��*2n!`n�����ݳ)�H�C���`�57٥][dK��I��p�]�3��}A��_Ѝ����CA���'�o�}8��{���SM��֡�	�3��y��܇�WI�]����
u�'�V
���U��@��9�z>�g�|�#C��b���Cg�2V~�
�W����s>�h��-�Hya�����j,����1�˅#o��6{\j�Oi}k�d���7{��wk���Q���-���W���.~�e���G��<H(����c� Q�����6׳�7�5g�Mrᗐ���)�ΚZa��VVr@�?h���]�V^eG����-s�8�m׀p��ܻwf�K���&��H���Q8h�2=���R��g�˰�n�%�)ei�0�	�Mk�g����^>m{ѧJi}�l~f��9�} t�o�<�7d(�A?�t%>��T'z��kk4�g�P4V.5L��jt��{�Y}Re����%p�D���v��a���S7F71ez�E��?�5��ԩ���,�@�����s��^��+�o�\E�38�H\����*4��T����]\4Z���(�W�݀��e@����zf�s��ɦ��r��s^ �=n��<H��T��>�C�]��ċf�����L����f�Lx�=@��F�䠌�j�ϣ��q}��f�_$�]c�.�]H ���}�G� �\���n����R���Ʒ�	��]}�[��w{��Q9�ܴ��u�ɼ�d�jAq�%I��H�)���L�Ύ�e=��c-����v�ԺTB�s7F���[Gߺ�G"��jUX�??*��f������G�i�8Ӄ�߄j��^��T{�pԝVUN��JP����C�R-�����6�@�h@�Uv���C�@Xٹ�1��4)g�q��q�Ƈ��4D1��)��}S|;L��S�9�%��Fd2P��d�lX�N�2J����W�CUuD�L�B{��0릳��*kN)�J����T�Na=/���q��g9O��D���؞�[^$�^����?طW�m> �O�#ӥ*`�4�8@ٌx��x�Rlz�T���W��w������9�,����M �x���<���I�ra+y]��8�,�hf��<�Io��K�0{#��H"��J��)��8m~qe�l(�gt�C@i e=X$�ּ��~-��%6��'��IQ�l���&�h�&6����@�a�Zɨ��)�h{�Q���k!/5�U�h�*>'i/��i���PΞ6��<��X�o��f	�j��x��`v��Qϝp�I�l�re�aݸ��,l�-��]�����YI�Myǟ��l߷7�!����ߠ�3��R�Te/��D=Fw���G���׊��?�71�U���dܿޞ�Yɇ���߃j�g2P����M���y\1���՜�&K�ϝ/�1�I���A�Y��� �?k���7?������sv�XkFL[j�8���H͗�r�L�{߹�܎Ԫ/��ą����C^-#��g��eC�暄#�xD��ӭ��63��5�Sj�����#/�~�ٯ�����D�yAm�8�WCV0�[P�)��2��= �њ�(��U��(�U�jX�t����"♍_�9q���1��_ź��/�|��җ�A��!�[D��\�W=&`<�Jƹ������U"0�����s�9�^�t��O�j��A�-W�@�WA�C�F9;��h
�9��Aw�5nb��q����-kL|s�F1���N��u��_ډ8=���*���N\nL�pZm�^����b%���wz��������l�,�e��{>2 2�q"|h�O��t.�8��>2����}��g�.��;�-�cX}�3��<�`ڞ����^��V-�M=���������u�lsai@�݆T�p�]�?�L�,f;}��q�G�H@�cx��'��1�M�=�il3�i ���4�>ȬG���37w鐜.̓Q΂��})6w^�B)<|��Ш�k�co�mD�<��:�����ix���-$�u��w-�m�|�6J�*�i+�����`;�G%����BH�â�IӋ�Ui5���[*�%���?pf���w�K�m�o�aijB��9�N!z�V��D���U�<���]����#?���>;2�����'�>̹��j�}bͼÇQ�g�y�I�ӬrIx�򠥛\@s��5��P����~���!w��1<�Q��ۧ�s��E��<�!էz������L�v�/�J�h��bHz��W^�ėO~"��-�x����}�z��)@hҎG�WU�WӬ5���T�
�t��a��LE�9\�z�K @+�!Wi����X&�uB�.�,�����^$-SpW�0���/��rN��G2�ʤX��M=`����I_K���P�,����ї�"��q�x;k%[������	/�{��}Br{d���a(�W{_R�oI�%p��Q�ha}����W<cF-��o�֖O\+���X�� ��L���;QD�?���r�R��~����n4J$>')m��ָ�
��"���R��z���t��|��"vYH�Y�q@��`͕9���a����}����L�B��02�t坧���E���%�;J��(�|n	�j���L��Ŀ�Q]<}�Q�_�g�9��"�L��ۗ�E�v�,�F#�e��a���.����]��̩�03]8|�є%;̈́��,Dl����)&{[=hҖ���|����3��nSƈ��ѐviqm~���6*Dw�#ˑ�uN���݊�Ѧ�>Xً�5�c�`n2N�����~��h�iO@�mo�~w�odӯ���w>IQ�faJL���N�MRw��8+Pwڽ#��������G� )�H�Lpɮ�p�].ݝ,A����]����E�+;ϋ\:k�z����7=��,�X��#���J�^�%Y���R���Ƈ�#�����w�f�I����%
	�+6{û�/h���.��f]w�r����۵��A��O�6y�,�V��}૭Uu��n��˃o���5Ɖre��>���@tJ/z&tkÛ<Q���ׂ6�r�g6L�[�p�t[��Q�![Kns�kSsy����Px�W��p{�E}���_�7�B�͛3�㚑G��zE, E�(�Ŗ할]qX8�&�Ś�C��oc�}������ƁC�̟3;��W��	W�����0XB^�+��Ha-�h�m����9��c��{�uǆm�Q��<P��mV9����a�U�d\Ha��K�'y͎����k���p�#�dѮ'�h�xS�����n�h7}�¾�_�����rX\���8縔\�{����iףyö˂��Wo�������BSE�\����y�d��Z�wt��:��HX�T������U�\k��j?��$J�t��������a��++@攒���CZ1��wd����ut�o��I�<���@f5�#��#{?D��RÞ�#�C��%'�-�l^7��M匡�����s_���y�$s�Ný�ll�!�vrsC�I�������ҦέE�.9ϩ!b��
R�Ҡ��G#��A����Y�|��s����UlT$�R�~�
Gx�
?���]^�}0�;�X�����&Clo��^s�Vd�91'[׽���B�7o����W�{[y(�nT_��Ơ[���p�a|3^AxlXׅٴ�}>�y1����z]N��j�@�4�3��ǂ�<�J�� ���:�5�Ҧ����Ш�[�&"J�z����!�	M?�=xKJo�C>��Q2�u̾�b�6�_�X���3��J^xoȎ�t�pużC�H�&m8�
mM��[;i}m���
k8R��'���zo"��Xv�h���VN����:9�K��%�|���ڛ��(�)��r6�`��W�-�8E+�_!6��gX0=�5EV�1�Ey�v��G:~��Kǵ*�TԞ��哸bDz��tBn��~�vwկ��1�Z�<�ʲB~�n��`|��Y$���%���=����}sF�NgA�?h��V�
�V߇�,L��f�|���t��̕����4!�s!��ȅ�<�d�Eڴ���PFO�׌�'Ǻ�i�YT�s#ji}lȯCV�+�n[|��'���
#+^,U�!8���
7T��3���./�?��\#�t��j�������;��,)���r�M��m̱��q�q��)�6I�#I[6�I:�=נq��۽+*$Յ��N�_�:G"�Zz�/��b��h����D�X�1Wۂ�1�<>�ї��7Y�=O�}���Ǌ��Ő��+�ߓ9�
O a��m�0Ye��Mwu�j\���t�%��,���?_�c�T�۵���m�1��������$��K�%�����g>r��ba�(q��,�U����u��w�?�le��I^�z%��y����q7��h�2��t�}9~S�}�!CT�ɳ-���M�j�^׎6|lg�wpj�4�(�R6�2)�֦q>>w�X}��OҰ��Z�S)��zT$l;�^��j��^*U��Jf3�,P��Ũ����euv�Ѹ�&�
�4�?�Q��Q�ub���G�g��q
�HN�������}���QoNg�����\�h��:.����#�$dbatn��3�j*D�(�O��uW0L�X�if<����8�g�n!��e, Y��o�b�j]����O�􈣮}=B��(8tj��j�b����$�Q�0�Y����\Ͽ<n�ɱW����P�W��O|�P���ycd7�݅sl,gk<E���4<���/IE��\bL��(�
h	$��+�v'�'�Cs�="������R2-5�G�n�M��Թda�͡�6R���ֺj	�6��z���C���%3i�n���&s���gN-�.���|MG�y������,�q[3�5t�q�G���4�LY�`H,�,�GV�u�Ů)�;?8b�^zMG��'�#�l���e1T�v�$�#K���������4�4����ʕ���Ԣ'�b�<=gr���>��l]�ܪW�ͥg�n��,.D��1$ ͪ��_��� 7��;��u��.U}mb!���#���'?�@cJ�u]�������A�<G��5H��N��Pv8�ܶ���c��'��֦D�?{nu�P ���^@��&�>�F���4�B\̊��.��.P��c��� �{����H]޲�E^�r_�(_ɝ7 ��5e�H������<�A���B`"�|���'J��K��yDӶ����Ӿ3�r{�r:��zP���w
Bq�v@L�����\����+b؎��?J���[�1붐�cv���[���[����Pq�Q#����fO`���I��ԡ�y)��Z�+n�C�������v�?�L�ӣ��cs��=���e9�$�o��3u���e�[�k�mb;�D�?��2�o��gcc91nv�Co$��/�L;��l
�z2uW~��߼Ƚ�nj���0�#���kM�@p�����덋�!D 0���@U$5iM���p�9����F&�(��|}���m����k�6-�|g��0nٓ��opl�ҏ y~H���)���X\����%z(݋��)D�z�����և����nw�b���⻿�!k	i�.��:��m��o x�I��-'���.�݅��M���mE19��IkL���=I������}���5?��zl݇������;[���?u CX�����FrN+}�K]�i��27�$X���@ ��u��:/w��C�)�)�M@�R7|o9 f?ݏ��;���p�`S��=�.x,ys�RQ´�c��sF�i�u�d��hm<&Y������Ë���y����޲C�����c�f+P6�*�nP������8���\�[�Ƕ����P��b�"n�T�̐&�h=��L�gk�%�녛�%������}�M(��}�H��A�IҴP�9ⴆ2t:�I\�hgXE�a�1�\��,��.�����@��qW+_)o	O������<"��C�G���=�|�W��� 1�I�A���W���<�Կ��G���3�k�q+�C�"$�\��}���q6��ƫ�2eZ������$U��������N�h��V��b���E��Q������;��œFW�8��7�"VkĂB����"u*��2C$`�f㉜������б�V�����>�gD��M��)�+��_�3}����,�PS�Q�t%W�
�J�����S�4�5�%4!2[4�/�H�7�����ך�bb��q�B,ح����W�41��: �@a�w�RW��M��Y���U`�K������O�sW5@�<g�ܴ߹��[��pm a'�O�ʗ�������[�����{}b��߄B��%�x�# ��[��ܢ�Q��|����A�M��C�KI�I���Eoi��Wc���@�	�	���A�Dw��F���(�)'kw��zD-�2B��r1�f�Ŗ[˔���ku�I�P\{��/�^㩮yׇ����m=�X�7�x|}��^v:��Y�=`�SeHP��~z~���2ғ�d�'6��b43���ڜVZzm�ߎA��lH���S���;�q�$A��LF���J�=���t���O�����! ��Ѱ���h��L ��[�s)�����viM p����ޖe�PKc{��T�p�%y��@hl��(�ʻ�%Ξ�uܩ�Bb��*�daR{ ����Y����ԽS�)'����a7=���qCu{�}�=L���f�g�	�����11��	�e�j�fGc�KöhA�*\~�k�#C��b�K_#�s|Yf��I�E���c.g��3���GօS���{HEi�16�UP�L��XV?Y��X���4����d67���hC�H��%!4����m�!D^�D�h��tA@/>� MW$�7'V���\w�?�N���}�70���բ��+�<��0yl^����W�I�*ګqu�b�^,%4�ᦕ��FKG��V��֭�d�we�>J*���5��Rɥ� �K����V�T�.�9Mf��hv4@m���w�ED���O*�l^7V����{(|�Bj�ܺzms��sT
�)��E�l�L�Q�A�b��F�[�l�,���EPx�>1��,�u	5$9��!�.+Qϲ6�Q���qΘ�L���-���*AU2y*�B흳<���] �C��~��1PANf�����O�ev�ϭe�����u�>�O�H�׿o����Z�� ��.$���s���a�P8����"A~� g��P��<�_�s"9u�Fupp[l�	io�z�d��'^�I�t[?�iw֯�*���AA�4��(G<5%�Uj�*|�P�������M_��wB�����^�?QbPy+I9g0=�\�����,b��E^'JP����ڽ��rĮ�n��]8��j�t�g�U���˂���{_���a T�%��Z��3��������ҕ��� ̻����٫B/���\���0��P�q���3��� ���Խ/6�UÎ�%�2` g盘�����L�D�z��Ǎ�D|k�m�Osc"z~D��,���M��5AU6^X0������@�r��!Ǉ=*d>�$��_}1��z!���b�[�e)2ۃ�h�F$D���th��ك~����������RE��
�,����ER�"�=�=׶��Z�((7�����ܰ^>̓�l��nAn�h�n'NJa�Z�M 9��(5�F}�Ġ�����I�Vbe5�J�v7'{�a|Y}+�S_�)�D��j2�p�F�åK�������������4 �4d�9������h�/!�!m�lp,R��{jR&�H�!3!w�f�:X�9�;R��~���>��:O#�|9�
�����z|�\,��8Q�L���m���3���tIQO�D���p^a��}<R�z�É�C|��
���w��G�t
��|�[���tN�6> �����j��&7��6��!��+����s?E���p��W:97�]��E�z
K���yc�X�C�l�e<j8~����b\�E���<eK�Q,�ȢO	����}��kٛ~+�ز{�O�삲M���� |@=]a[���C�vleޗ%�~�*"ZK�*����R7  8�kR�|�Y��ʯ���Dc��ʰ��|F6�$[>]����l�:D�,�u� �4���ll�	�I!z�M�@�d��`(aY�=1��A�PT8�*(k�^�V�W �
H�T���8뭝�M_��Mz��|C�[�ʶ�֒Ĩ��g!;�7�;�WY>Uc**��+o�
�w�[�n�lΝ�|�]�Ѽ���34A0���5�����}��3�ZQ�OY5��ˮ�����9��f�
�V
V?Y|ZB��LE�pCR�4y\�E�3�/�N~&�%2.���UW͢Nf��"(~ ;�0��-x�q��
Қ1R�z�ix�pܡ������c�%�C��!Pf�Ӣ��v�̭[� ��������zD�;潄C�MP��uleB�7�E��/u�u�I vh�<v�hL�������
������\���և��b1bE�ۭ�F��<E���o�14y������Y4j]���QTN+N�Ya�߰�6A@�odRְ�I�� Pa:��)�x��6����&D�} ��	E����}�:}��gn��M�tQ�J]�T���������qq�i�� �e���Y�4]�U��,T��R�R�F"�Ʉ�ܐ�_�8��y��GyF�	� ���* X�ᴣ.�c[{o�g���E��]��܌տ7/�9��X�V�l�,ѭZ�ף���EKyP�ۺ��2�����-�[T�f�M�O�:�V}�{���i��������7�-���r<��|�&W^@��d��BC��U���!�֚��ؘ��I�n�S���ɺC_��8��QlT�,TT�ڃ��zG���\ֲ)J��1����J�v���'i!�9�l�c>or�X൛�6����MU^��A���dW�QE���3e�3S�n ��	N6�� n�(ġ�G��{��_J��8+�<D
AY��/�
�na\�Z�e{���?N'�#��<~��//p��Vp/�y��:5������ὴ�8��EM%z���j��\� w��t�6��J�PD�Ҽ�B鯱gYφ ��M{���q��Z.���b�V��(��ڷ��Ӭ�6��hh���=U"�f*,���6����O�I~����?��<���_�	�h�[d�wb;�D��J	������u5��P��M��w�~m~A^C�NQe��,s��^T�?�Ǣ����o�x�1c
�����Zw�a�hk�q����Q�=Ӿ�U�v�LB���������i��<N�2�ô�-m��_m=�!�l���x2�Iqbv��20}�b6s�yƺ�y�w�u{�;���<q��eP�a�~I۪?w^=W�������Y�Q�H�In@r��-��|&���~2�l��4'ws�}�t�p;�'V�0)H`�@Fޘ�6�{u��-X,����6��$��
����>��鷋0h�G��T��_��°݆�E�n\a� ����Mt����Gڥ�;@M
{�f�f!�M�q��}w�f<��@0�u��7�����Ow�A�p�l���tDC; �i���Wڃ�%{29 ��{�� p��)9%��N����c,�
��B
L_]�0�6Ӆ����y�,"��OR�)]dn�ǬY�����5�i!?Dʾ��+: ��Y�� ���!�.��珢��6�����"ڗ;שs4��	��}YO_����4��!�"p/]��AW̺!Q8�����DWD�$3�}� ���%���t���E'��#}`��\���;��-��l.ˮU%���R���	B6���c��;�ڊ{H��IXЬ(�Ӽ���.3VM�v�&��I*��4��OO���+�9u��F�2�J/��!/�����n� I(�f@��i�'�j�Hw���y�A���C7V��*���YU�>����=��=>��AM�� p���e�ݮ�͒��ڔ>��;�BFBH,Җ�>E������%�����}+���M%�*X{^��OJ��`(�tu=��e���tW6���}$J�(�܁� dm5����	Z��	�����e[Մ?O�r���
��(�X��\��zH��?D=����O��zg��� <��Fj	�O�|�"G½HK�>�`�9�Ib���^9�]�^�ih�/d�F�q�ۏ�n�JL��uK�1���ʦ��b���Ni������EƫOZ<�����F"ό��p�]b���%����K���K���]�{�ƣ�U\�u=��1���K*��N]J)3	e]���ruƌs���s߸F��[���R2e[��äV�۔���;D۪�6@�)g�X��8�w�R2R�g��4t&N^UyJ�{ZBQW�*���K��5�}s�+�AS+��a	R5J��%e���D�݂ΈR����F���i��&l�d��z+Ñ�&�M89�9�e4�{(#�.	A�w���R�
TM-TU��T�6��_��k�K}9�/:f1�l�J�
�K�a�_�a3P��`g�A����W�s)��4`E�K�ܒ��ӭ����ɝ��97�
?I"�ԙ�(��R�v�����a)<�\��m㭗-ꋘR�έf���Z�wN-jo��PiD����f?�tGd+,�]Fm�"�C�W�ȹq��?�#��r��yu
���M��%���-y���gN����2��;7�u+;ݏ���C�)����W��,��.G���Y��a)��Mg-�ǌ9s�e�ˮ�x��p���3�����4+ݮ�F�>�N���wN�VFrY�Ԗ �MO�G>�lWm���� �� �f��?Y\�$��#�;��^��Jբ��	�O&�V
�7�R�O�	����E|̯i�z#hN莨ߍ�l]��ޜ���'��5�-����C@¶#%� �:�AVF��b�&+���w�y����҉�52�0:R���/�dX$�P4X�P�`x�6�z���ɮ!�U��L��_m=��I��!�Lym?\�ǂt��#]3�J���	��*y�3K�~���r@.>�'�>��k���k[��O�gȗp�O�)r�d������K/�j*�Y��|�����N����|^ʑ�#�.(�.G��Sc�L��r�`��3ZE�{�3T��_~'C�#�'���A��g559���-����Cֶ�7;��h� �v�� c��b���a�:ؒn	{�m��?�=<<��v=�V��d"ԩ�$������p�0��ɣdr1r���?d����		#D�G����wr��a�f�3ϝ�y�I6J���o�����U�'�I&�?4.>�&�4����7r��{nÊ�}��,�a�Z�� R�Kڨ0�����n��{u�#�j�D:8���Q-Y�z/���sz5%��i�+Y�Dh��oKJ����Sz�D�1{��/x��r��b�%�C�V��-�p?�,�F��!�߶II�e�=�߹���
xg��/-��Иl���N�����ɡd���s��kUx��PS2��7��h��?<�t�)}f�!��8�6g�5*���i'�n\}|Nvr2!��?s��h�C��������xv�z�WP�`}⪩���[>��b[�Q��+>WU���2��t��{&/T^�KsR�$P�n���X�>2d�_j��Xʴ�����̡ȳw�ېV��T���	��۞ԉF��ɅO_��X�?�$��mTR��Θ|����Uv"i|�pb:/����t�C�ϕΜ�T���	Ee��	���r��-� �/��E ���M�D�GϱwOՅ�N�l^�#`EZy�I��:)y�R�o'uy�;�N_��b$��r6dS����ۢ<6�O�X��2�7R���ρ��������J�ss����!qH��6>U�ɷ��%F6�-vR��X�*�t�*�0��Q0%�D=������.P�����^�w�*��2�
*�e9�1���2��%2�)sW*}�����Ry�5�T���7����m�%Ӷ9�v�����̉7Be����N3�S��F<M���F�%Y	1�Ł�LYO���;ysȢuק���Y�R�CyN[���oFy(ֻ�Ԕ�<���
,��[���滐3XF3�5nfe��F]qZ>/ {V�?��T��,yy'p�Y�����L��d_�D����K�?��l�3T�xDj�锕�L-��E�?��<�V>ן��m�ԭ�k�qZ�D����
's������;�[m2�;s�a[b/||��
D�4�^�����yˤ���_�yW�"k���PB{����ͺ�hXϴ���*�FU"|��oR~����~68ՂZ����i)t�7��f���~�T��<�����}�	�X�i��ÏvE����7K���idmo���⬪fKd]ѭ����Tmm���|�E��?�����ҏ���'�Y"��Z�w�\�1�����Y�]�d�e�xB�;�^խ9
��D����7!�O�d9���4�j��u��9���oŖgk�fXh�KrV(R�߾�F%"��JԸ���0����N�TF�����,�;.%�=`�����3y��j�X9ʮT.E2�%%�����q)�@�K���|].��^�
z=̋�KA���J�/�S���C
�@��m^�hm �h~+�_�s�!�ؖ��P�MQW�oY�Y�/J|��\�/4�hx&,�E;�����*҃[)��c�\��0�����z��\S�������?KE�ī�	ʮ��ؙ���K�.o:�}2� 
��#�}�2OutN�BW�%�������;[�Z�U�o��k���j�"�� o������<�X�r�����wF�Z4V���[��á�q�ؕ�-4�tJ�;+�؄(���$B�~��Nm�Gct������መ��h�r~pLM�`M%6.K:��X���F#Yn�lXkx�D�����nn�r`�+C��9{�.@C7��*���LKQ-�yԙIc��(�y�w�y�~���1��Ē#��b`�c�tc���>���Ѣ�A5��g���JH������ٟ�>��jM��(N�$���lu����	�K��u:�-{X-OjE��pbၩ�ce_N[������9�"vk�,y�i"AQ6r�����2-W�j��F�J�l��W	��?DN�Z�?5Y
R��/���ʪ����u�"���
RuJ¼�"ʔ�
��H��:�-wZ����1�<�Q���M!�b�"w铸~�Z�.��ߞ��/���ѷ����*���gk?��61���.>�~��K>�^�|���WB"'��RWi5��i	&i��)yDCHEWH�K9��7��ȫ�<��V�h�q��]M�G(�!�����7Ϩ�3��Fz��
�(	.|�~���c��Y�m��{ܷ`F�?��z�B� �z	Mb31x��s5��*Oc�|�sK��@��WR~Ց���|ߙ��I;*�ܮ�$��/�>�s'��*����-�^���G��m�J�-�}�����t�*�n�����v��i����ɥ���V�_o�J���pR�\v0CMQ�x��%&9&n��:���c�X}4�*��!������_Ӿ�Y䜡��jR�62O7õ� `�M���Ε�e+��vj���2�����^�{�b�uR��e�n-$�&��-�
�?t$XVf�C�k�K�+�G;�fpm<�e��Q��{9͈�"k􂬸j���ްu�1�F\]p_N��rF��q*�.�r�Y��.�s��`e\kՋH�{7P[.�V��ԁE������C�k[tYa=b�s���T��ﲵ�:�|���}+���/�e�'숷V-K�5o�`ظ�W��XK��F͙<9��H�{�?Ru�@2�x,��{�T����Y�b�!�J�ǃ���uֻ;���OKWv�ss�sd��-_�����$!��m��S�;��������Dpmg�\ĵu�]�{�ח����Ù�*�V�s߿{ԕ�:J[a�Q����!_��V�+�οE�8����E@q��n�g����\U�����&�Oо.;}��Ʊ�m}���o���gv�O;�y��9fW���W�X/�bu!={�{���H#-�3�e׹��ø�+B���U��~K�\E��u�s:�Y�'e��s�I�a=2d�"����0K�i� ��q�.˪ i��-R�O{�'o�y��^x˜٭y�O�_g]I_��z�b�+:Z�;hy�'m"�g��FD��+ьؽ��I��O��Mw/�J��
|-����5l���yI�����tӖ-����Z��T���aI�f`��g_tt�N2�̾�ZSƎ�?�	Yt��z/�Qe>��b��٦w8���C͙�[�-��n�Oz�	���X�C$SD��A;��_��.�̬lX���L��)<$���f�,���t�/�;j_�}7f��߲}���9����W�`��|ΡEu�S/� �`��c�U��A�bQ>��6�-���-B�z�o�Pʇ����+g�w8�o�7��<G����?�a�E�ĵ����Yҗ�%�+'QM;��ʣ]׸���ԣ�2���(/FX]�R*�zf�,���G�Z��sn���'B����V�>�搴O�/+3����%I'�w/�ED�L}�.�y�Q��=��||�8���jFcqE�܃MS�>IJk�����̫����
��FL�"��vS�V̺�r�-
���3�KD��Y�.m>c�`ZCM���X�� ωΫ�yb!bC}��!�յ��8�켏�H(��4���Y�=���pV_�zee�7�l*x
WB���@(���?����s���o���B��5/e��:rժ�˖�n`��e����&���^C˼��5��rϕĹؤ�Ï��?�j���[v���w�_�6���F&�্�E��rT����h�zZ�0a��=���n�i�ڪ���Kx���O��l��皅�%��3�5����������`��s��A[��X�	c�e1�9.��
�/��E��J�����`�v%!�}�L�Q�]�B��r�6������Uw������Q��hΛ<LB�{��GG+
��(Úә<Cm��j��=�7Fe�������j��Ml����s���H�,�,ɚt^����aQ�]ۃ���-*H+
H+ݠt�]*�94 �5Hw%C*��94�ߞ�}��x�����^׊s��\�x|�b-԰�7P�SK��ju3V�_�D��v�ǭoB�{��ů��c����Y�.Z�7�!���F�j����d��r��~����Hq�򑸸���&�f��u]����m#jN�Is5��S��R�7��L>�O�����w�Y_�2nF�q��/|#��]�K�!�+H����ڎO�-�����H"���ϗ^������Lx_�|ҥ�2��������`�l��
����Ս$>`������|��q�Bcu԰���]/�{�،�BG��$�Ƅ*�8���eH!�ז��q1�+��8F��z������'�w�F*��"I�9D���M'i��)e̤��Hܣ*J �֥�}�o����������l�����N\�1�ARnPM�}p��Ҁ���I��|�B`,#�8��<!j	`�g��
e1df ���J�N\����Ё�o����ZP��=,�Z�B,6� ��,��G��>2��&�F�t�Z�֚5�ҥ��M�ZUl4v�������j��k�$�8�H!�a�iޭGg�R�x������+�}��fedj�mF��u��|�rq�7�J�9܄c8)���u0�.i�"�<}fM#��C|� -��e#r�)��[������Su�g��n�o��N�d��R�R�jX�Xgg�0҅w�g�^{�����wi�5�{Z�־��EѪ}��0g0�l([��|g�EG���u���l\)�ʑ�:��r��'�qQ�	nM����{���IsW���B{+��ܞ�J�K�Ano����2�Fʐ9���f�! .�3w������,)�1v56U^گ	^'���Wx��c�w���=��U�dy�k�]R�y!C(>�C?71���c4vP�t��{�����c��m�������	a��&�O+h��T^.2_{�;��j���&|	���C���m������֬�U������s�=>i}�^��J�������)(X�P��r)�@}]����X�y':7�lP�ܬ4���"3h/ꖂw�Jx_/R�x��2R4�%���
BC��p�D_CP�aG[�!t'ld��,vס�4��z�߄E�'��Tc��1�CW#B��@j���N���zM��M��ff6={3�O���V�ޮ1�;@��]�QU�q_�#i�M,(����?��o>K���B��ۨ�&�"q��e�x��:�H6��z2&��&����(@㦚���i�z��A�Q��b?�8����_Rɡ�"��Ź��wXك���#T�2IEU"��s?���V����@B�9X��Iˬz�%T�� �c��i�Q��Re�x�˃�v];�@t�i*��\�tU6ͮ���5�����Q����������� qe�{�'��vh�?�W*[i�z�v�~$��j�� �_#�#=�33:ȵ�W�'�i��:�j����@]sL��Mm���4�:�ڢ�(J�$n±|>/�,�"��J�!�}(lt�w�1ԛ�F���7��=�n�xY��K�5�c(��YŒ��ٛR�� ��G��P�r!����O�v}���2a���y0����� *����Y�ڐ�i��$����Ħ�p���U�Y <v�x`�D�Y@�nJ�Չ"��8l��G�	�$�]]SVR��DmP#�q� #�˖_��r�@�+uM���2�Q�44��LH���G�6��Q0Ϩ�L�B.ĝ��ߍ�b��X���s!��`���Kp�e)�Cz�l�̸�˫^��dVz�r���!$�#$�����k5���E�`���>��1���|��G���i�П��I��j�%k�ʁh�x *�:�����Bü�U��������l{�h��xf�hޒPtfY�3vEh�="Wo���a�:׆����Zl9����8�>�J�Z��m�[�r�����TY@���Db6ʳ*��(�R��	\�u�4�K�ƳHV2�t� �E8�Z�uT��B˟�~ҟ��7HC��7���~A��.�2�$��F��Ifw`��k���h��+��1���ˮ�cD�ܝ��)�Dt0y~�v/�k=�,.y���}�B�����\�k�I:s���X4S�����z�/��	�-�?�.�?����%�6��
T2�%�'�4���J����o����`3=�y�yC'K�o'�����߮��P��/#�Ɩ�,R�M6W��)���'\��rԠ?=��%r�ɱ~�_?��v���qބ;6�&��w׀�G�t;��~�Ѭ7 u.���EHv��i�S˫����=^!�[�v$6����^�_:N �1�����]O���Ҙ��I�)g���/�HxI���ѩlg&��ǐ������~r�/ɂ���Ҷ��\Dd��c���<~L��
�0G8+N"K��W��$"~f����Ђ�/7"��D��l]�I�a�L��s�f��Ǝ�����xJ��!I�N�=�}aCA��q�ǥi[�R&�U�0!�"���~� p�ب<���
����ir�	�p!G�N1����6��{��!����R�&����ˉ��۰��G��F���15�##��|�з��m�� P\��R-�`ܞ���?�Y�1���eV��T��
׽�ODp7i$��q��AΦL�tM��Cz���H܍�n�"��c�鹦{vcD�̥�0a]+� �M 7�3sXX>����s
�����qoX����,��S�]B@���p8-�9���:���xo�s�F�{bK�g6@�p'��Ў�.>��?��$8�ё��F���B$N�P�·���o�v�f���]����:�U��ݞ���C�K��ε�!V������Q��<�w�G��q���{J� ��i�%�M��Z�j>�4X:ow�b��/X�CP�?ӟ���o����M1�������������{����;�#W�*w�3��x>��3��� x�&����a����/��Z��9׌�%�=�1"��H��|�u�S`�ߠ�!>�X�wQzSw9Dۧ��{��5$q6y:���\wA����we� �.��٥��/�~+�FP����-�j�Nfr����:��Lp�q�1*�ώ	�o��Q��&1m�i��~��eW?�����0#��jA��%�oU�N�� ��}��k�9k��g�ט?����Y@��k(.+v���I�i�Ƕ���DA2@�� ���4��E.
H����G|s@�{��9�eG�\����	�3kT�L}��XW4�na9����;���8��:a����զOVN
0x0S���@�xU�oTFX�6�Ȅs�Uq����'=)�Ɔ����=c8��pH�u�� W.���^�\��Ƨ�ILW����\�H���es��Wpx_�@4�R���
dJb�\�������IVp�p?�ְ&@��Y6Kj(���6g��	�b۟�>���X��L� �nf)���v���6��[����lY�x�k�3G.ɦ\�=�࣭�Ll?�� K�͢
��I�m}���?r�NT
�S0s�̳}�����8*��HRQ�نl�]k�mJ�Q� ���w<��7��������ɋ*�<y���[&k�gE�g�ɇ[{�	u;
�D5�]��:'�� �t�Q5�ʇ�O��P�+��Wr��;�]�T*cD�li��X�)�۟'�����a�.Qnt��Â{ѕc�7q��KO����`�;�]��Ӟ�����28ٟB������w��15�+�)b���@qLZ��ION����)���Y̈��l�~�m�
6��+��s�f(<Ȑ_`F�:PbG�q�;ޭ��Ii�(���x0 F
��� S���]A	��	R/ `��{������]'0���02ՆIzV��vS�\����	{.j�*����dP�P���JK%\h�������r��M�3�oH����J;�$�C5 �o?:��2��<�e֙������sk^gk���w挞?�n����������e�bb��1
��^ m�?�"���ۙE��D- ��l�{Y�2phx���eL!c<P&�>�����G�� #����F0��}&[!���hl5 �v�F�,:z��]��}�kNem���}�MM�9���L�؛�cJE����������v���������gM7��Y�%����W�k�,E�H�e5j�x���
6?��ߥ^Ti�������V�F�հz�|���I=�Z�4b�&� k��&<r]ߥ�����й��	@F��+Ϧ}�Հ$�C#�F���l΍��Cr�pS[78j���5a��οh����� T�.䯶SS�ƨ�/f'1jb+����0���Sz�հ�?�Z@����{��J�Ȓ+�H\��O��엢X�V���KPK�#���rޑ� �qW�����6���F�����\�Y]����,G��C-���#"5@����Z`�*D y�r|v��^�S�o�	�ΫO��N��B% ;<�@�p���j,��Y!���{�����1�1�/����V�*��m�Ll^l����_�n��m&��5'X��>c�ܤ�G�h�W����"�XW�Z#Z� ��?Ru#~?��9���!"�y�ra2���i;|�;ke���S�	$:c���]��̡��|���whAB��{��ƆLH^��K:0k���P�����m����3}8��%y3� �[|��_�3|!��]�hi4V��Lɟ���a�v��$n�]Ǧ�+d�\�Y��W�y\�����|Q-~/F�%��n�������ˀP_�Ϲ-��M���-]^��Y�'v���~>f�r�j�BpG!5��.�-JX�t�����S�>�$U��s]z��{�V��gd�
,EJu���m�	I�w��xD0�MB�������M������&\g�\�]��r�I�O��~=���/����A��.E���L+�Wa��E��(n��m�4���|��gυ�e�)�M������"&����z4 �d���$�?��sn���<��uX�T�q)'�o�<!�Ax|��^T�h��l9�j�������y��M�~����mn=�����ϲRf0s`���NW���ށ���|�`�R ��xz�\�8���	z�c��kI@;r��<��[���ܕ_-�
�M����A���[��**`�=��YA�W�@2�aي��,p���Xp�
§��k�x� ��=�YE���o�Ub���,�}�*W�*�)>#r�rP|.���\����`�V���e���o����ԑ��f���V.:��B��mǡ�q[E� ��E���\�������{\�q�~Rȳxr�f-���|̍v4͑?��	)@.[*�e'�%�8*��Yrs�K��)�͐��3x9���*�HF����:�Jc�"ru��r6�V���{�'s~��+��43�&0���l�㔠{і&����wҢ���˶��l�;p�l�~n(���JZ��%.��-�*b��d�Z�ڣ�!��J@UJV�]7v���+{��xEY�4�*�K�}9u��B�Z�^y�̋ �'��a�$����a��}EN��粦{6C8k�����	�v�m镔����O�,D_T躘ϊ�\�)Ff�k�6�v���H��g��� :�M����D��]s�MN�!>:�*5���`Z�xW��;�У��u���I��Utѣazn/���u(>q�kl��:;M"��q�=	X���{i��qw'կ�����-:�q�痁�E'k�M��QGEq�t�<_�`J3��5	j_�>-�]t%��F`Z�~̱4Kh� ��V�Ǿ��e�ƾ3�ݱ�¸�y=������t��5���:�|��s�5Ҏ��ڢ�5���.)Ώ�nӭS����j��A::܇�|��?~������4�S�K�Te��Ib�������o1[�|:ox���/��Q�]��ʾT,����N��}������~7�U��ؓo���N��
1���~~�uL\J@e�������}/dr�'��b����������]��ޮp�_5����б�{���a|\���n�g��h��G��+��f�;S�3�grL�#��<�&P]?�?���y�����)V�ⷺ�q�|x���������2�С|�Rw�ϤS��Ej�N�?�S}�.7ڲBp��̦�Hr��?�^�	���Rjm�HBUeͶ��O��p7i.��A?���<���x���a߅���9ѓ��}�RS����W�G�:Y����J��&���0��%(�{i���Բ;��בrQ��d~���G�ү�Zat�!�4����dH�+Ԕb�>s�U���o-#Y]��{-�7�8	J]���I��F�[�1��6���l���Z���45�*X�^��9���F�"G��/��o�ѹ��f�3yBY�|���mMJ'x)�H�`f�ڿ��Tdsl0y��͉�߸��w4�F�蚉��͆?��uHb@^��e�Q ��W�5b�l��Pj��0�"���p�˗҃Y|rcϕ�4~Ue�: qDk��_MLT��UlQg�˼%u��~����lh�gs���K���^��/	�@�s�˘C����D���볥k}��	=��GH��ҪOU�$�T?��g3U�F��-[�l�ت5��vc��,�6b?�5��l�F��c�(֥=��ЦZس��;2�ˣK�{�<�S��*���쫍���x�
���-o���ENW�2���J���jI�^��Kϡɫ�����?�y7q8�%���B'1�,��M��%:��CU>C�=U1K^��j�<k(r�(p+����d5?ey�\d��Q��
kO��s3����q�|6��ٺqREk���zĕ��cj)�A�y6��[��n�1��#�o�=e�,���y�kf��`������!0�%l�|�};�p3y'bG��roD>�a )ʦh
�݅]���σQ�!���i:��p3U&z����}��4�+u��XuT4RV#|=����I ��[����l|�I,`z�T$�����*�q���ע{���bL�I��b��p�Hͭ���c+�^�b��X"X}���G�)<�����iI�L�.�3h17��c�ehR��������;6S�_���Y�M7�*{�#��������P����=M�87N͔[1�l���͍��fe�"G����fމ"��tQ�G���f܇ѩbsI�j��LȬ��ٝ��-k$�����d��e1�Vh=R����#M�o\�\�d���7��l{��&t��4���ury�x�r�ޮQ�T���Ǫu��4����Q��p�����X�1[�!�T�E0��_��F$hvk�k-𲀧�*��]MsOi������m��<�VZ�Y*Z�3ü&*�����b�jɦ�0dUQu5�#�)�{Y��/I���T�o2;9ޖio�����)w�W�]4{'����g�To;���|j�#Xe�Z�ؖ���Z#�M����r��֖kw	�U+n'��vw��=�J6O�Ƀ�wqXn��V�M'4e�\�9LO�
��ּZ<�1�[��N��st�⇒gJ��.&P@�j�=>J>�1W�~c�}j1��we
[�m\|f��B�-�߶�r��$��K�����^���x}��E�����2eP��F��z�r�0���^��d��N��{ޡ��5iS���W�jk�J0��6���T�~�r!�67k�Ko�C���~��@�ƴ��>��`Eb7`
9�aH�ܯ��:a�7:RC\��/��u����%멡�Pf��F������j��>U�h7��n�ݿ� h84��
.4F���c� ��cuI����]Z��V�n��靼wő�P����^�����;���T6M�n�E�x1��Y�S����{�!97�}�&d�Ƒ'S�*�#Q��X�:���2ļ)ɞ��O^� Uyf�`:N�Т]c��C�ՙiژ�7�p�UD*��M_����l:杤���#�"�_�#�o��F��7.��zU��
4ׯ�{�/Ja��TfX%��f��wG
��
��խ'N�g��7Om�o3�x�j�F���0�9��H+����9�}Up�{�� `�s��X�BT���5������3�Dq�Q�����v���8���c�p��������}����=������m��󪼸'JUc�qo�Y(���w)�3yœ̜f?����6��`��A�H�!I�4��j1��ؠ=P��g�+[O�$�3>eX6�ux�f��Y0�P� uZ���Z�,@u��['��)ļl���l��k׊o@�1�,�u���Ň(���WN���s<JnZIe(-�/���C�K,����S��Ν�����h��N?\v��s*{���m�uf]7+�{���!^R8]@���O�Bc(���������!�1�S(��^L��/s�?NK<�<�@��޷��q�'��Ƨ&LO��.�B�j�`������v�
^Jֳ�K����8��Ӣ^�|��F�r�	��80�+9�cN��q���.�-}Z����R0Ꝭvo��o��G�()3ʵ:uv	�����#Y��}�U�V��}�Tɲ4c���x2�n�'R}��5?�U<��X� 5��W���*�_-
w�ލ �Ǿ�{w����Z�y)VI�����*|� Yk��G��y����;m��"շ��t��e�^�^w2�Ui=�>ڞG����u+��U���6��2~���*�W�"�ni��ѱ�����	8�	N��������	M��G��W��±H�^��v�hsh��[^�M�ӗ_�8Jє+u��e����3 B���o;,��� ���V�O�����
�
.�ގ���-wL�=�qx�?���J����+��^V��H��/N�x){m���U�S�]�-u�u��=:��@��t���0����A���M#9�C(Z�ka����=��7��ڝ���S��˸��6i�}ƇZ0��%3olH|��58�Wz��䄥#sX��ͺkq0?ւ<.D5k����+�ā�7\�Bx���(fn����WN[W[y����n���%�!9$Yϻӿ�q�7pn3_�x�]��jlȵl��[�$��'��c74(1Gl���|j�U�mt'fzn�mf�?š5�q�������U���gU�ܭ����R�g���k�VQ�{�5[85�mX��}H�9G��TB9\)8�B�r �߹�S��;��o@�i�Ywg^�ƾ !-;!ޣ�Q�d�����
�fm��Y��_�sm	��K^�7��6�*#��U�6M�C��xu����Z�9'?v	"u��R��V�0(��25~�itUm;k?�|���2W"f���oP7���a����z��#�#8!�����L��ϊ�[�"�	7<j'M���"}Y�)0.�_'�O����z�5ea(.���l��R��V����9�J��g\Ay�|vl�u����.�ݯ�U�k"�C�{�,H��ߚrP�C�k��kl��2���ޛ�
>x\~-e\o�'�p�݄�>���*�y���]әh8�w4^U�&�p��S�H��m[I2�t>�lw6�t���uD��[����������:n3*���#X�ب�?W����R�������Y��f�˛�>��cu��cqt͛�����ԳC��s��x1-z�}*�P�K
U���4���i6�Ǻʄ�=���]C�%GAȱ�&)ȕ�<��� �i�T����@H��>5"]�	��[`)-�I�1>�	.$�̱Ǉ��C�ŭ�Mg2(O-'�O߬��6�d�N7Kj��;�YE���C,��_�E}���Hb��=`rF%����+�����nsL�:��N1����E����ً�q��I�[OԽ]tXm�O�RS7[�3���p�L�?+��;�&|�X!��fJf �U��ix��f�M��2���/�i#H�4�qA���"��&���d�{;Һ2d�b,�=WID��Ĉn��K�����)bxJ�+�9�e,�P!Ӵ��o��/����w��l�x�y��ӬXagو&_I��C47L��v|#.�,��ay5�;�hpK~.:�Ԗ�N,��u�-�QV�\+3Lq����a�:�ӆ����5T3\g�k��>��q���7��`�8^9`���*[�f����~Uکg�O�p���_G��sC�_M��<�E��,6�t/��=ߢꝿU�;1���z��)d:ڬO6_���3��G�W���5=�q�f-�Il���!�Yn�6�LХ��j�l�	i�4���i���X/]'|����Й��H�O��J�����+��ݏ�����%����zކ]�t_�&Ԇ���4IYW�B�].� p�t�@�7@��ʴрU/�A�-#�:���VoB�r&ZO���9x�����x��*��F��e��z��)NŠ7�<��r�@��m��.�g8n����z+5�^���̾�k�A}p�p� Iw��1����~��v<���*�7��<{��Eŋ��@�^n"�/-5r�Y�}Y���W�h3�3 L�"*�Fn����'�:��9H�u����Rbx�_�|�g�цm������/e�d7�:�F���^�6C�Y|P����M��䆁��>�����y�Bud��{�M��05TJ�4�dp�!po�����-�Pe`v��z���ۄ����0[��(�����R�(#A���r����cH���j���K<��l��GėR��:��Tᓣ)eoҡ6�9���I����[k&��^��x��U3����%��gQ����ns� �s��(�S�s/�����K��a���.���|�����G�z��RDN��:s/�!y8r�WW�0��б���n�1',�輺������/�+���Q���Ț�Ιqe��_]�;"�;�V�<@�� =.�QQ,��g�!�2�1�yu�[�+�|l���;?6�E��.��s|�.�
����!�A����'�d[�����|$��=��CH��\�	�����[���Jg��!y[O���٢�H��_7_�VC��i\�d�ԔWz�
�����d�|�r�3�y�FJwl�.��D�E�����h��l��h�S�B7�>L~h�[?ᷟ8̙��-�.���ۏ�D��e�uҧ����=���q��P �B��X�v����hn�5P
W����Z&Y��n|���n���^��R�e;�P5�c^��եB�g.!�=�
5�y��^���(�B�8��k�(^��_���D�g���Ck�͵le�W����ս��T͔ �iȉr���T	�Y|�=
4^��F��y�O�0m��b�oq �$�f��w�!��x�4��͵��mZzO;��gF��5�
V{�.�6��+�V�a����|���{ϑb����x鷱}\�w�y��ק<UY~�J�I{; �-&>:��cLv.~�+�����+E
�0ś��p����|"�k��%cjX��a�n����U�ӋQ�[��{˪%�z�}G6��A6�����;�]a�ٌ��)8���Щ���R+��3��~�i����������r���כ�����;4� �"s{F��<;T"ŋk������=�sU�g�Ha��	�a�=�i0��@?������V\�m3�mV@b�b��Z��أ�|�����g�����E��<�O+y���j.�vi�B_��r8ד�#��s�ԇ�
��6H�䏞����p�t>���` �(Z)����2�@!��yle�C����VϷu���ک;����1&_W�.E�p�/ae���3�Uu���bX�Yt�'���+�p�-˪�����1�L�Sp��zq�ucm~��9�0���uɄ���fH����/����`���7�s������.=�;'mi��Ƀ��5�H}��Dh֨�uY]������MMP�zޑj����طN]�Ң�D�K������i��t�����ks����|�]�N>�v�+��y�î�r�1.�!��P���� q����V��B-�
vvG�#��
�:p�f�M
쫄�����Z�?�LLS&�;�00`�w��8V(m��*"� �ʪ3
����q_-%�x$��G|~5��>&�o��d�Ad8Ya� 7:�)�����/u��N�{)�]��W7���Hf�`Jk�L��#����G��̜#��D���r������:��<���wy�L3�Ïv�g���ԝ�s���5��`�7VZ�
gu<ť��y��(��1�7��-�D��Ԥn}�<5����ob�7�$�k*b�����AYo�8bi�T$��v�m@����l~F�w:5A�.R���:JqP��$�v7F#\�9�l��H"zN[����$��}�DN��5a���^�p��{���+��}��?�آ`�A��*��{e:ϯ��f�ݥB}O�|+�1]�C��A�k�(�������ŗuf�t����q��%�ɢ�9,H��0�';�+���F碹@u?Hi�+���M"c�*{w��_�s�Iq�,uLWL�o.�H������}���D��W #���!��I�U����Q�1ý��9;�E�%�_�/�d�����
u))��;+ص>(ay��z`�WVV3F}�k����5A#?���j�"���?|x�C_RXh��P۰��ț�๛���ǚ_��cA1�����K��lWJB���u�˾�)�K����qN� xOÀ"�k�?��C`��7LK�&6�:oK�W���m�����6Ԁ�]՜�T�V�4e��k�)Q8���w|#F���o���f��n��>��O'bdԬ
�YƩ�������6�m���y��Nan�@Rm�*[��2c9��d�gUw�1�N:a�Ȃ<xn�č�9G���)�������˪���$Fw��ߘL�h�-�d����?�y�4>�Xz�f�>S`���z	z�C����Xv�3�M,?Ğf��k��~��g4ط)��ˌo�����-|1Q+��<�������Z#2�P���d?�})vY�fa7]o���n����1��E�y>|I(HCl�����k�0!��G%�h���^Q)�v��ۦ:�
�!���5��k�f{J�,�tr8���(W��H���f��>^u�y�����F��0 �9�2o �8��_V�]��g�*���M
8�.���\�ۯ88C��?�Qf����#�3K\�/B��44bc���7��-K��%G��Sg�ݲ�-�8mp;h��TӞ^�}���h��i�عu�(7��cn;m��Ѝ�y]��()k'��Ω�%$�,]�C�Ƶ��_��X]�?�3�)�+����mg1���a��KY?�����ɮNŮw���^-��<8�0�?�zu9�X����yo=_i6:Qw<��d�����4Y֣���������*��ܬ(�Xj
P�t#KG��A�	�-�`,
^IR��J���'�~u��4�R0���&��u`À���'2L�8k_���lʻU�Y����n:�v*Y�W�S�K�K<��7$o�(4���<z�XA�x������[�W�e���s+˚�P��Ǹ��kQ~QE���;e�=!�'��a��͓�ҡ��#��y��ja�ȑ׸�p����~��x��i~��{��ce��说��I�U6[E,c�󾶺� л�:y�洛cߋ&���d�.T4@B�Ȁ�Ы�{�kg�I	6�@/�n����$��1)ְ�P�����A-��%k�V#��LSg�139�ku��SR�*��w�.s��p������\�$2�ZU���~B��ɌQ�N>�	r�x�_��υ���=�*\�oO�S|~�@	_��^�P�߈̮��q�u�~A=�o�\�@'������wY�cOk�#����ꎐ9Qb�QZ>#V7�>��^�i?���HrT,_?ț�W��z`������\o��l�j�7ab��w�If����w��&����d��7Nji)�$%�u4�߷���N57�{�-���׋�z�2�x�D����45�J&�f>m5�Q,�K�;�b��_h��Ƹv����vU6��Ć�>���Ԫĥ�^�aS��G^�B����`����ʺKq�C+�e���o=4��6�/�2�_�U�=jӯ^�-�r޵�����0��ۖ �p����w'8�IqZ>�����o��)�Q����xcQT_��#��k���뎓{ݷ�6�tB���{���Vs\V�{�NV(cO&����5�	F0��	�i�7�I���~N:�J`��<�2�?���?��������^�n��te�F�[��:��<����e7�gS�S0�¤]#��t%wu*�}��M��,�Y8�ߜ�We���a[�a�ȃp̃Q���ͨ�1��w���됀�^�+L��Hl��5,Fb8�2Q��A[��_x|Պ�.ʔ�i�
0�UKH:����^�l:�=6���W4����t.텕ӮO|K�UF���3u��rp�ح2Pzͷ�5x��A����ubI��RR��!�TV��CCS�9}$}���	��*���>
��c�R5(8��% �h��Y�K�SNov�����҉y�n�X$erK���-"��.�1�n�8���=8�ߎR�m�(t���
���=�Dk�w���#F9\7�D�!Q�=?� �;�4� �b1�TfƱaQ�|J��~�ZN~Q���18�^C��a+
�E,��0�cI6��<b5a��z���t_>�^V�CwYݻ:~? �2�z�R̼L}��VL��liD���=��J�q7)�k���(�eЇ(���|�E�BȧC�.2��s�ï���.zqB���D��E�����U�mԠI�=}�,��Yfү��A׏D1��/^3����0���G�8��nr�~
N�H������LGǠU�N׮�'S�`Р���8k��Fk�X��f�Dú֣���ũ8�T���e�������nY���B���Tw63P��S�X:��X5(���Z*���-���(l�v��b���e�t��L2�6�?��{��7�9�9.q���׻���3��#98��7깅��|�S>�9*޳�&e��z�6jA�K&@O�^w0AT��IPA��S��^�����\c��w����
%�EE<E��b����ɫ*���gC3����uRuQ�e蘯ʬB�����r���Q�F<�G�\�B�,���w,R���gS�k�{�1��'c¡ڔIɡe�NB}� ��kS����F�"�vh����h%F�����Ļ�-��<E��*?���ґF�/�� �p`�8�<D1$Uq�@@��qz�LF/��J��� ��B�D��ܬ�R��{��@ςv�KƲ�J��03Sõ����4g��2���;���=���=�r�\-��;ւ������_�HE���7p#F9�mݩA�����{[h������6#_�;gP�.�G�o=�Z ~�a�{~Pc��I�r��<��"���jk�~u��Q#!�9l16ȣ��I���;�*���WqX|��v�n�j��Z�p�D>�Q6N�o�
XK/�`���Z	f||$g�tx�$�9��� z&d4 :�H}#����ǭ²���T���Y�~����ɠp�gE
�����ޛ��Sݳ�l�%wF��.������b�貚��u�oK�ϖ�D'�=z�������J��m#y�B/�6��Q�"�\���r\��70�OP��Ҭ6�X_��^�g���:�_q��s�_R�2�p'/�F�I�=���Ai�{�0�"0c�����bH��Y(�l�7�K9�t1��=h��	t;�;�«)��Fa��=���iF�cmT�QN����%~��m��/#��x�Y��眝�s �/��x������č�e���e7~�x�ܶ�~����-h�uqp��<;�R��|��6豓;�P/I*��n�[����{�g��_����r[Ͷ��~�Ty̯ሪ��9��r��깾
��0.N�9��7����q1#K�.�ت��ݓL4lR��} q�����[.�i|$��<������'X,�mu��'���c�4ru�2mTƄF���S��(�E��^���J��J��B!��`������Gπ��3�M-��)� ��m)���j"�g�^X�s��w����(Hb74����i��w�a���U��ԉf�<�
�E$��1�i�����]�t��6�ݛ�_�.�s�9�d&�w�=���а�\��2!�A0��o?c|g�ډhMɷ�~��7bD�}2H�v�tv�l��<1�d�f;�<a�	�R@��8o��|�|�S� ��˝�}�tQ}��/aZI���{�&�x��eUT��?�O"M���*ل@� �����;�|UڰbL�����|I��;Z���+ ��E���_�P�d���Ė�Ie}u�}ʩ�c<Ps1#�����PO����o���cp��i3������&�ā�C�vm������W���I�%$<�YQ)ö�y)�Z��8l�}�2�R�T�h�*cXQ�M�@cq�����x�*��
����$����e�frO�KP�p�{����r���P�B3E`e�~	���pP���<���/�I�U"�ܷf;��@ͅ�!�dƐE�Ҹַ]�6�u�޳��PfS�[�H�T��T§gʭ��E	2`�&kX����sAIo��!1 P��F!�+�d��J��xc��氯m��7 �d��M�}{:{@���oB�[XZ�Uƽ0̅�6<e�\9?� ��H=_�{ �_/E6���a�����i�ͷb5(S�����qQt�ۃ� �%
�� �JJ7�"�,)a"!)ݵ����HIw� K7,������~>���s��}]���!-�9Źq!֚��F���Q�y���i�Y�e�j��-����HhI�IPS�`�����6Ԕ�Xy�	ւYR�z���ɼ�<^����s�i�4�˦�#�fV�TS�@�<�W�&c�`M�@"%�t&&���`Zsǯ� F�NN��������+֫r�VO��(|P�&SJb�|j����B����w `�K�e]&{L��%��dD�������/bU ��8(W��vN� �\��W��r��U��M��?�64�3"j�^,x�m���II�T��@5_	�����Ë���9Q����h�\�z��l@�B��#�L1��\һ��/�X1�Ӕ������g�%�����"Rw�V]����	���� fI[���ج�È�w��Óא�ߪ�
�����i���sɧx7� c�-��6F3]YK�/�G�1n�K@M22HOX�)�%��N���Q�8���seD'Q��ڇ��U�`�ϰ�t�u��CO��ʫ���@��ʟ٣�C��UV��Ǹ�h&��"sF�S���o�)��K	8r!x6��8$�ڂd	�ͥ��k7�����Ɛ��g�4	�_��?��q�Y�ɳ�1:����kyB!R��P�=|���-~��ܻC̥��!0^M�H��v+�xաX��l�ZI�v$S7�;P(	�WA�'^���g�>��	�"K<ݤ$��Eo�Y`��uͲ��;q��'��8�ix�dW���O��=�$�u�����ń�Γz<� _�\\�sU�O�m� ~��X/����e��9{�]ѯ�CU�п�S�Yzt���o��7U�W��b{�,�%1_������dI��zP��_���·6�Pg
h,{w��·W�(�:�5LP����W�2��ۤz}K��B��'�xi�< �46�K�9�}����7�U��Fzŗ�<�7ƫ�	,S��u�g���9���{0��XA��u�ax����
��K	q`쓊�sgDWn�D3J�|4�����J�?��{����)oM��չ��Ե�$$μ��7��R������k���o"��a0�F!v'hK�n�� z­.=I��@��7d� ��&7���6��f0�8j19���v{cV�����J���o�9ʍ�m��Qa��g�h�s�X�S�.H&>!ǷnN�C!���̈́� �G���Ҩ]�q�8�˗���T��x���Qcum��]%��F�ü��ݢl؀DF�X��{�Q�\��m�6�!��Ө�aD�zLf��I�|�:-TbLf�K�Eh�pD ��(��h�l��� ���?w�b�1_�M���s�l0�lb����ߣ�{F7ΙQ�ǣ�=o����(+	�X!��n��G�z`m�r�i
0��aH�v%1�H��JȊ�˟I��- �����7��k^+�}�~��Z�����-s����%{�t�MlLI�ƹ��C�<.�d��P�?��=4�!Ubm!�X4H���Eא��Wn婉�/�
��B M�5������@���Q��:�,��$�s���xHH�V��w��k��ZI�f�@Cqݤ�`HDEY��h�U�~���Y�3rfEw��x�G�)�.]
����F�7D��|1��q@�&�(��jAI+��R��V�č�%C�3���ş�� PKU��	��3�*H���^[Х4�`�R����ȧ�:���~S�������|��2�������6�MQ�t̱v�r<�j�����N�04G��\�gf�&�����:���7 �y�eR/Z$/���L���j%M�1��4�cl���v�{���
��"uxs�����
��g� d��`Y��m[��7 �|�/�J�@]M��R��[k] K8/����OH4OiiY��aϿioO�9%,�M���y��Pkz���tY8�S%,3�}yF\���E�]r����|)'&�h�g��]V����v�Gq$�B� �h՘zp�:�&T��'�庯��4ӝ��l�܎����>����r�냥�r9OG&���[;���b�@h��r���6��7l�N|���z|�h�#$�.ԓ�F?쳸vvU�_K&�������_
�ye�$��X
�r�w!�p��3=-��
Y<�u��/> ����><g�F��A���>�O�sNCB��h5�7�A�ԲC0��"��3�+�q���|H
���ѽ��=I�ck�+��``F���+ r|Dv��\?��fd�����Z� (��fp��?F��k���>�'W�ƭ6�-�,���n	H����çUU^6���6ȝ`ǫ����8����֋�fR��!���R6MY���(�:ӝ�ֵI�-~�^�Ec(fN��c�W��{��)�<&��Y{���F7�s�-��0�4���m[���a��ĝ���9��)��2�Tn���>�Zs
(�T�������� [�A�j�%B� Y.�Ӓ��qa ��H��P��v�%_)�K:d#�A����}��j��)�-��3���_��Fʻl����8���`������w�I�U��Ψ�)~9� ��i�.����?T���P��ԃ�����`@�����N��T�s�"ϡ�ְv�yc�0�!Z�hX4qՀD���,&����i~d��5�̯w$���:��:�� nϵ������l��Z����%X��X��w�B���F�4+���s˒�ͅ5|����⯬|�����?�\���ֿP�{&����b��@n0O���g7� ��<�'6ɞ�� �Rg��P~o��Ng$H����Pk�K�h�0~�0�T��gҲ����弒����W<m�x�?�4➿��\ʑ�ؤ�ƫ���h�ǈ	d�$M3�=g8i8Dww+�-
�`�D1i�ʋ��c�)C�HO*��]�C�~��>��$�u�~[
��/䄐I/*:�6J�:��(k�d3��P�� ALxD7"68�s�x$-S
�U��ȃh��eU���Ld:���.�5S�J5�L�hQmyzL�5��~D~.���,�/�k���6%U�.���橨!�,�o[��8�8aec��i �3N#�7]O� ��F�9q�D�>��έ��	h�_j�z�H�:�^�E�$�G�\���)��߄[� ��-y^��O�R5��^�7Ib	���u���bZ��n�7�����)|��d$��](���Y�0x(���4Xc����Yp�
���cNd?���{���?E�?� o�j��~�9/����s��kU����B��q2�,�PzÃ�A����H(��P� o$���8��z�9��{W�Cx>n��d�P�$G���+���/n����Ȃjz��1\�%�ɛ�1l���q��7
Y�u��K��O �'��kK\�h�*���Au[^e�����򡋏�qTI60#���Q��&4�@��h�A���|�?F� h��%v�������q`ԋLd��\a&�e8EV��W���X��&�7�5��)*���a�bpo��b��S�>�a@�_1��&ʛ����Ow��`�ÿ�ͬ䉒��E+�����d�Vt��k�L�)KY�����K�7�
��h3��` �����fv���QkmXǙ$B�����0F���C�|}�^��~�oߚ#ܯv+����Җ�AnB|���L�L�*G����h�G�ַ�YZd_.W�dlԓ�?�'` A~�ʒ}��E
�H�B	N.�[ pN��U��,*3�������:;<�(�>��P��F��5�:@e(��Dv��N����m���6v�c�BI	��T���h��H��Fens��s����S<ؐ
��o�~���N��4���t�1VO
H˗o?|�D�vU|��q�:���c�%��5�1�l�7��~d��@��־�����k^�6���!>ѽ��e�z8�%w�!9b���R�� �����kÎ>�0A�>_��?�`G���7p�(��52u�$n�~�-n�]2
�ND�����̸�p���,Vq�>��bae���b)X25	!<p�
S3J�e	^%�������x�ziD�o��*�����x��y�OP	�=���6���>��C�4>��	~��j�I��/q��Ӟ5�g���ro��yVu�Vt\z�& ��c����u�r�����
�A�:ncg`)�Zr_m/����Ƚ�G�t���~H��X*m��o'�@㿉����~��m�z����A��<NQ�Z=}P�U�s���;S�k�шLq���P0|�z��s��Uh��P�ac~�_~Γл�ZY��P*�e� �\�>n� -�FP
{���Z5?X�7J*�Өf<EPB�_�(��@��`����TS�P��%�	H\$����h@����6�q�ă �ϡ���4��������O,4#߂�������A�b�z�A ��g�x �^8�8�돜y����ޝ/�B�r�'�oui&�P�觥�)�K����3�����kk���4nL�-��H#�L��&PǕ�F�P"\�ǅ,ZA�t�Ø���0Cm���c�N��ѫjSPہ�����;��U�ux�΃Y���-�.y�K|Gw �Bɨҙ�|E��v	L�R?�;h9Y-�b��v~:��#���^��u{�w��	Ȝ}�`�[�rp_��Ǟ��B;�'p/Y[ФG8��HT�I���_�v{��qeB�A��"t������D�.`!��l!jg�������j腎C�'����n�4�c��I���x�j�D ���lp/x[}R7���.z�֝������ʐUD���<k��>Ðp*%�����p��Bkr�ZO����7�^�ϳUO
��}[��i#;h�{�F��͇Z��0��}@�1��	�Z����H!������ ��"훓@V{���f�*�w���C�E��$&p/0�X@JY���9���Y�Sk^�_�,]ĮL4���jbՐ�5���Ӳ������í���Z�g��|� G}>ힼ9� ,�S��E���r �K�6�r윑�hD�`uˏڠ �`��R���oM�mC��m��fR��{h��1�A���p2��x���M�w>}@;u�{!6�8z&�{�gn�j�G�u_��^�����1ho ��k7H)��)�Q���<Y�m��QI �Y%��~ő1\�E#vڷM#n��
�'�mS�Z�v�j8а F�jh��f=�=�ƍvEV��ނȥP���K��ܵ^�+Q^mmn'g�N!�;��>��9��C�DQ�P0HPF�ê3��KM�m0�Zn�Dռ�hr|��)�8 �
6�b=�2b)y���R&�ò��ے���'>5���4�7R�o�JEq��2x8�b�-��r)F��n&��@��x`IdjF�v�9�$���d��Df47�q`�n�اhgvw�1�*d?�x��Zൠ�!'3{Ug�ě��ຕ[�3y��l����:fY��ц��Q^��_�'�:E&=�sF=$ގ�˅��0�gn;��0b�1$��<]ᒻ�&6h`�у��c���ב�C��k��U��?o�8bޢ��T�!��"=~�;����0� `�3P2��}G�
�)�gߢx �
�
�5t�t�����[�����_M����>��x��á��ò,�OG�3-�������5�𒾗}<�����ʹ�-q��ԃ�{�\��F�#I��]���0p�W:tn׃0����N��X c�W���z�g*pt! vg�y>�Q�v{1K?�hH���L0u������W�W.����r�Pm���vKtH�F�:L0L�"�ky�6���(�g*߁jٯ!�@Vz��P�֚�e�]�����V6��-�ЌȪỻ�%�r���:fAtޞ���%�*��B�cS��1p� +O��xq]��S���EUF1�h�^d�� ?��bm:�燹#}t~��Lr��[�}���򔰞'_�Y�y�	��*��f�B<&%X�t��*��'�#��Z,�� ��e/���}�����w��g(6��1��\˼P�(�Ĥ�٬ M�_Îf�2�Ə�oJ�|0�^�g�}�d�%k8��ih��p)��t?*T���C�U�{+��Z2s�	{�F2�ȶA��@e�7X[_��mB���m���M6�@B����:/$\�C�������]����la6e��X{��I	CM�����_����������ti�[�=�Cek���T��wx��w��l]�kS�{��#�\ ���h��^�Yt�`��%8�!���M��Rێ��R�ZS�����b�y�n���r�e���{���������iǶ�)��Ǻ@�m�[Ww��li�����mt�v����B�X���������aWQ�M�!qo�$w>�Z֯{ծ��Gz`0��` R^ğ��D�������6��c��Pl��;�l��j����TE�mJPS��W�-��Vy�Hm;�ؾ	�,��Wc��Ni[�aP������&%�\��^�꺻����vLץ�|R� ��$|�]���������$s�-&��#��Տ%��J���]��E�6@2]*oaS�l����Z7ASV՝e��m��~ɯ�r�j"ɨ������r��i��p<p��J�k9�k�F�_U��xņm)	
��pcC���}׷}�I����@���ı@0�c���;�]�$ʮ�"�S��Ed�Osɘ5�	�tf�櫛�ۃA��	m�����u�&,�6�ի����<Z�~/��~�D@�ژ!�k�)i;�7^�rWp%�S�މb-"�+������JN�?yΦ�Qc5�����j�y)����폓8����Ӆ�|D�Ӻ��Z� D��y,/l�86A�|o'^�.|�=��D]�JVW4�Y��إ՞}�N;��}!dY�0*>�8��ۺpwl�����du�Q�G�J �.��q�Q�ʙ�_��ٍ����a�Q �6�S�=�v���M(�k%z���:���:�|P}`�!ɩ���Y:
`�0�!��/��<.�ٿ[q*�����
�.��R���O�5^�ҿq�h�<}�y�-c�3A7s�Щ](
�X
,���`¼,v����RϴK�/�]}
�^�7�Ć�N�]/7:�f����s����=��]ʂ�@"�o�<>�_g�8������[�A�v��w ����J����&	+|�cR��F������Y�{/�A�z)��~6�'y�b���4�?Dq����}�r��5���c�+���u���_C�D�3x��0�6�����V������a���vM�4���q����g�_*l�ksJ$;%����
@ZY�o�jxR
�[�2F9V����k~ :0���(�E�������,"͕W$��^D��;��2S�7징�ƴ��T0j3��GV{Í����o�-�����(*�%�\i�%;e:>c���H����>�4���Y�J(y:��T%�k���l��I�8"H=�p_��3���WӾWx�fQͥ4�n^*vqY�`�]u�+7}���t�]+��9��b�Ҝl��0�Z��{E��~��'�J�{�:�{�P�8�i4��o'�t�˓�w���Ffw��Y
���������#�Q>�C�4�Kcb%`<�ґ t!�?�������6��P�'�s�' �f͕���
/Ӹ������2����.�u#^���ɴ����p�O�s�[vj4�o^pH�p��Ps>\���~!���:�=�7���o����,����3\wĊl]��+�&uzh��Z��� �P����k�عoG�օ u��^Ԙu���ZF��PR´�O{Z�b!2D�"�HD����ꉮ���~�벉)�ub��XN��׻N^�����3����翯bcb��ÄU�(E�ػA�W]����?�m�ΎW��sMM~�5l<����.��w���T-}^�N��I;%�x�FN"&���w�{q;i�Ck+�\9P���o��LƑl��a<O$=�A�G�Kf?Y7�N[s�VvYg���{}I�ȡ8������i��%;x��ktq����U$�@��qR5N4�_��0���Td+�=��ʪ���D#rH6�U���q�'ve)�Sl�tI���}�}]{��6aK�����2���Ogoqş�Or'[�T��
��b���G�}�o�!A��{��'=2��s��������kL�/hw'��N�3]G�s�̞�7<\�$eP�hr��;&��>r��^�.l��V��O{�+
Qtk"�� !��i�K�����=�w�$��5Z'rF���w���!�8Wĳ��u{�rq������oq���1��B���ڂFM�/*�(��)��㬢9�hr�)VgX��{�Z���ǰ�Z�����8��Q�9�1u����Mǃ.9�+���Z�YiZ�-HUA+�k��f^u�$��V��D�������﷋Mݦ��7)�3c?F'�/&����'+E*S!|�#S��ĽmL�����'�����]ы[��z�����!��\��ϥ���E&������1��e�~E�����ʨ�JYE��+����`�s��]�����ܼ�5?�M��"U��	"E����B57 �]2S$�������R�OKW)�|L����*O�O���{���z�}�Dfo�P��Z��ؠ��h�S���N�q�ˋ��ϒ���J�.�*�q�'2����9�U'�)R���Wgm]���PE�
��Y��k=�Ǻ'� �B��{1u�z�&:�ؖ*
�8���)\�z���[}����W>��h��M�ʦ��i9Y�ͅrm���OM|
�lk�W��ck#e,"|]��f>z�R�no�z{\��:�P�63�w��$�a�rN�c�{}f �GW��8- ��v&����
�_b���T��k�5�\�7GG��h*�'��X��Y��*`f�Y��搉��HW<�Wzz8px�^�Ơ#���:�k�6⁲!۸r��g�0��� ���cփC۷=��)���L�� ��Ϣ�-X՚�2燄%���A#���<�����6)CRk[�)���?Z�nN˚�E���憓p����d_��$ke�WK�������L��w}�Y�S���ʗ.�o'��I4=T*�)H3�#.R�(����9S5ߤfH0�7]�箧X��˧��Yp.B"�ܭ4��7�F0�O)Yz9��_ zr�{���������B������!"�x�K�k^��F��D����2>�~��ge�"�ە��浢��ւ^[�c=�X�U;3S����K;I�����V�
�K1LH/�})7�ہ:6�J��h� DH(�6s�i��;�>++k������1VUQyp�|�f�%{-s�X!�,�82g��:)�^����@�y�HHC�ߑ�zu��u�Ae{�胼`#�^t��YŨ$Ի
Ԩr��	U�����gc�?�\�F-AV�C��]�b�_��SfYJT-��d,���BA{�e�Rr��:8��X�4^Pޥ:&�[f��gy�6��YP�Ց9�w �ʱ�b�Z�/�@CϨ��l�բ�4^W���Zh�U^Tn���kՑK�%K��9�?K�j �v��o����kU?�Z����G�c�G]��UvEr�����ϟ 6z��&<�9��^�Xh���4��Ͻ���EA�f�ٔ���Y"7�DezV
��R�k�T�*y�U)��n��\�����-t��=���l�}�)Sja)�z���烆����G��)�3Qz�*�3l<����L�[As%`��8��R���?0$2��$!��:�N��j?�H�j�6D��l\������./��4������:��8��K���T�\��Z#�DpN=gÃ�G��S
��f�+��x�+���?�Z|�	H�5˦���q�wϛPR��)�M2�{	?|����{!�百e�Q5|;e�H
7����d��8'I���|��k�Q.$��g����S�?�0��5b3����P�>bjI���p�~��8�����9� ��n�[�zYsQ��S�	3��5�z�
��M�{��&�0�"�S�9Ę��D��PJ�.��"�# ���Q+t�y�/p#,R�26Ϊ�pe-s��_�>���zFD�0�9	ѝ���".nzCO8D �4j�aJ��ߞ۔�.�-M���N%3	R���я��+�Y�}c�sK:�)��Wŉ��I�z@��� ����a^Ǉ?�06�f���0��6nQ-<���g>���R^j�q��`p$��r�d��W񁍰W?�(�X�7^� ��kq�1�EGH�B��.z3�.�ŷ��ĳ���U��L�B]�;J3;4��@��pWXn\���O��wM@mV��B��4\h�ta�5�#�]���x/VkJwێ���rⰵF}!`JŨj|K$x5!j�m�kC־��x����"�X���h�焝]|��?�c�ٶknz� �~^�������k�c���U�y��ٷ�E↢&�+n+/���@H�8�E�f���,7m^��������Pڱ�1=�#{� �l��kk������U��Pl���N�YجU��d_z�U�n��C~���8�M�&ƺD�u�[E;x�o���\�EÎ���&o[��(���� Z�����H(�'4����:;��Cz�wl�F)�
�mڼ�xl=*[��d)e/Ta�7/V��+IՁYY�\�`5"0�ɟ�� ��+v��[)�k'':���oKg��#��6���k��M�)MuB�/�e�o}�bϥk>�c��Kc@m6x���<昜r�wݤ�U�g��݂q�@I-��6�����\�չ��Y�U�B��'�I��肑GU��oG]��c��K����M���y�6��{6������5��K xc�6ǋI�{����}b�C_m�][4lA�4nt2�y"�ٛ��Ȁ�cӕ�SV��Q���M��Gz�й��f�v�"tw��纱"0�@W؅S·��i��f��4��^���	ѵ�;D~a=��y�����Ŧ�d-��h�K�C�>[������U����zh�D8�"�1�i\��XM:�
a"rւ�AI\��c���-���1ƫC��k�s�=?��Q�S4k�Z�����k�'	���|iԨW�N{z~
�-q�9e����~9�$`�1|%� 4t��fڷ�N�ϟ�[eg����g��f�����e�Z��7�$���f�r[ts�m�����!D��	Ԥ�:��ڷȗ�B�	�H�ӥ����+���rK�L�i��tz�\�m��GQx���_�_�R����2�&�]~\L��]����_��6�`�VHE9|xK��5h�~pB�r0_� ޶].����p���Y~09��X-w|.�����>l�M��
NktR�b������uά�����WA�������Uћ�g����#�֗�mM��ra"�!Z?���)��Tʡj���<w�s4.7�i�dI�2��,�^3%p)�Y��E�G��Z��G�ᵤ����`O�BfJ�z��`���+ů�\�--R�R7?��p�����r�~@N��3S�W|vڎP4�/�]�.?.�Ӈ�R;�a�H��?�%9�������U`_���uʴ���6��BPF �x���c^�l����?�\�)ձn�0��gX���8��y�}�Zi@��>r��ō4��)�y���
e Gm,P.�b��¶���&Fxh"�,曽���35����P��7���J����W�~��R�E���Tu�n�y_���̟�xѱ�W-��v[��ܘ��s�GZH�p��C���ٚ�qW��I0��H���A��W#?��%l�
'��&딍X��ISZ�7�?�:#J���|�Fr���J����r/<�pѵ@��l�s��UͯM�Mt��Ԕ�O
��1n�-��ؔD���b��=^`%j�2��^�M[���.{��vmk'c!u�ꔤ��O�N7t^�
:(��b6#�1���**ۙx;���!p���V��.�|������B�e��j�u�M��2Vf��E�)u�d,v���w⺙-�V��;�p�^�rxDn8>>��
����akjG�m�?Q��}���o�����v��D����M�q]�%O.{y���u5_�3b�K�8D%�}%LT+�D��${K띃K}�&�%�W�L��BQ�N���XN�ח�̕�7p�뀠�j��Shm��%�����؍GεAӗQ���΍oM%����5��iJ�"P�I9+�\_p#�D''
M*��atj>�e�s�;[��!E�'�\8�L�[��+��R��_��
�F=�SU���:��t�W�7h�	�����bA�έվʯ6nt�k����>��5�TNC6d��O��Lm��|*�j�
�����/�iČd�'~��M�O�%l��Ew���wvnR	�F/N�<�%S�viKbc�}.�Dֹ�!y����8q��ݲ����`���jͻ�S拕*���#��}O� zC��>É!l"	X=�^C3��9���3�!K� �V)��}���=���8�Cf�K�غWm���Hɛ��� ���J@1g*����LU�МzjT��$�=Ev֞�U��H-�b=�,Ǜ�!�������go%a�:�ʧ�ş<͠WlR|�FO�����|$���*'n��#%�"����D��}L.*�L�v�݊��.v�c��O�����X��ݚ�y.CY��D!|���2/Q�˽|�[o�H�j��/M�[��&�Iu7�̯,N��+�;���3�̕L��U-�D	;��H��%������Ζ�E_=O಄ ��Pq>��e�<6A7���p�pas�y�-ݺRb�Ӂ����l#�m4�O���2ꈸ2�G��;^��o�q�aS�E�:XI�I�&��:�WEg���1o45�(QY����zLa���,5Ә�E0s�����A�7Xho�ܚ]�<��̇��Gv0;��.�]�8�':�8��=�a�_M&�-���_y����P�ss"�+��>�BI��0��V#\|˩GW����ja�q�EZ�U�㘔)��"���;zgq����:Z��X�X1GE'���N� �FEk�/SM#�$�G�߉:REy�'������a��Nb]�M���*]�:�jҡ�/�%����;F�61�x�VZI������,��L�,�iX�<N���V�s��f#�6�; P���T[����	�)H���x�"P�gS?a�y�ǭ���nr���u%8�W5K_�)��h�D�f�W��7��'%a����uG��1�W�T���8(���~�餋����
,^�濒c)��1�MAF��̓lxV�ă����.��J w�l�����Z{&�8?�ؓ��}�n-))�\��^��4~��
<�I:ߙ�'�n �bno9�6Y���˖��tcپ�-!ΌNvҿ5vSSP
�~檿�8�P�C*�tй�_���Ͷ�����/��X��EWQϣ��D�9���ŵV��=��Ro�߫�ZT��j'���ά��;������|j-���g5V�*�S���VR>�����4�J�<�m�g��%�[5ι���!�����_*�2�c���l^u��t�j:%����Z[�.<cƮV���Xݫ)�V���>t�fK���L9���S�J�#�EmL������T�o5�������<\;�����9.轁pUZ\/�������~i�\O[��T���2���	�����
�a�)�ƆZ{C(%L(\�~�G���Ĉ���ߧk�b5�Ν6Y�~��rG=������P��Pbt���G��[�v/�\}�q���{�mb����"��V	v�I�S��i"��x��I�-��	�`�G�v㦾���#���k���`�=�ٔ���#���[�f���������~lɶ~c,\��1�[�u�H�"���v�RH ��@�K��rܿ�� Xo�	̷F��v�>ipn.���y��u:�����?G���覵�3���2��I�� 
釂xCS#�]���l�io�	\x98�Sm��h"���S��^.�ۆ���dc�>�|b4� g#'�2���M�q:k_�о�XLeA�����uyW����+>5Ϻ�343m�����ov�nsv6���Q�1Y\�!l�>�X<O� �� �@��X[�-�&��Y�$�} b����`A�'�=P����������݈󆧍�9�E��iM��.Y�I|��}N"r
Awbp�=����;�������O�Os�T�֫_�f�&c��f��%=����	W�NC��k|&pb�Gb5m��%΂��N}����L}��-P�����O�_�1T���k�`8�l�egz�vz��Ru����뎎mf�k����3&螓q ������Y���&�Q%�J��i�cq6,�7A4�_��l�����O��V(�_� ty��71�`��ó/?���@Ʋ�����������sT���`B��H��{}���ʴ�sA���$�"	`m	F��?�Gz��ېj,^�!����Zn��l]�T����nV��G���|6���.�1�#=ui�=���S[-ec����h�2�G!}3�G϶kS�5s��Mw�	�r�=�(��ܖ��0�����╌��}=�WI(�_~��|�b�u�δC�5h��{^�R$5�K/��oՄ��������&č�8.�:4-1.4\�}���3��g����]L8f�L`=��P˄�3a�L��7>��+��ڝ.��M�߅������k�Bd�;���ż5�}�>�`���� ���M�!zq��ztX�!]wǩ*�x7�J��U%������~��sWO�M�f"#U��C��U�:��h�=\bذ[/�����|����{ff�>iZ>�s�UyW���?7/�3�/�7 *����n8�U[q�9��oZ}6�%ηQY�G����!������J��j� c�qPv���T	_�zF�
2X�^�c�Y�7ٰ�!R�(�N��΀��ٲo5���q��vCߎx=�YŶ��i�MB��ym����~�Q��n�ӕ�,�Q� _��eBWl����L[ݔ�]������6���b���wW�Z�
�J�K��:|��t:��J��+`\EN��[L]*���vA�]�Q���e�1X����y�1��l=���)�p!�7��SE��I;H���Ƣ�;�T�T�8a{�Б!�7�f�R�ʷ�a��%uСńm�����j��u�XO5ԩ1����68 g���Mg
~PB"��Z�̟��H�A�A�����T�̐+�r)(p����dϜb�j�l�����ݶ/�t�p�峬V��O� ���V�����B5<��X�5��Z�:�e(h�i�rI%� PǄ@z�od�����N/~��{���~Y�����ʲ#�%����zD�ӟ.v�=��U%�x��wߔ<����z�i��v�+�5�'�ۯ���l�Q���sI�����M��"�b� ��M���.Q޵�˳��w�u�W��=�0�:�_GjtSL���I�Y��SF|<�2�H��h`s'�Z|?]f��o�����X�̘ޗ�)���!�����"���b���]��X#�Kf~��Z/3�S~�G����b3�Si���~�p��$��i���O�j�}/s��Xt�C���ؕ]��|��ǗV/��ocP�7���Ik�*�xG��S;���9�,�H:6�t�O�*Vܿ��iWJ��)d������n�i+7(x����>����Ӳ�x�Ԡ��֨�)l����;".�7[�/��7%7�ۺ�y����<Yߪޅo���y�7Z&�c�}�CW>���h'c]��rź�RbdT��J���C��z��鶝�`���,�U�e�Tb7�Z���c� ��i@#(��f�ӏ�/f��S}u+F�$�����3���ː�w��~�Ǳ�ZN�[��o�7�EY���۾$-�PJ1X����q8��n����ka��C�4�H�d�o.2�Z�`R�_ˠ 1X�1��A��W��D�>�ue�`a��`m���e�xR���#�_�/l��xC�c��m�6��I��/������,D�	d����]���5�}�����i*�H��S>����4��B�z��^��q����~�ؔ�8<~����[φ<��iB���m�+�),sc�dLե����uQ�9�8�;�P�l���Ŝ!��~�t%�8�����%��^�<�Ϙ�z���!4Ҽk��-���D�x+�}����Д���9�"qY���9�@
��<U���>n��`�A��֨�~Fqn[[p�@��-����Q��nn�me>������g���_G��6#n�������r� )��Md����9827w7�@�}]�1S���	'G��e��BwX���Œq�]��e����%���0�V+�ǥ�4B��o��K��P�c�7�`ش�����3r��{�ߟ��������Yf��J���ħtl���0�P�v��7⾡��"���w�m`-���YYuD�7{�x͌0���g<�g?�"O�M�|��O��K�'@���S��yp��K6Q�^;r:��l��.���h�W�$朠�F.�b/����t�1}\Z5�
��Ð_&��fsRGzD���>�Ҽ��#�@.��u���v%�gI�ƛ�_ e�����R��ɢ]������r�I�y���B�e̟WU�i�Hl���\�����^noWU�,i�v��Iąi�1�WW�����T}��Qr!���׏�4B�N�Ib�֥��]fwB�NĽ/�������^R�	f���Yy�X��?|�O+S��1b��?��y���3}�~�]�6^<(Er+D���{h�J�KFJ�v~�v��W��� ��`�'��)4+��F>������"	�r�VV�j�S� ���u<��c�N��R~bb(4��.�X�gHj]�f�~��en��[۴��'sx�ç��-�h"�B�C��:��������4�A����]���kC��ǐ,F��u�aU�_� "H7@��n)�i�n%��;9t���[��A�����������3����k���Qn�n��������W� �<�K;��,��$h��еh�T,��Oሟ�2-�큯��-ꟹ}���nѨ�0����E��Tx��`D��-����r�C�6t�-�r�����-��m� �&u���u,�W��_0�bc�g�۫��9�=	f�6[�$-ILM����b�x#q���"悘f�rh��- �@לfúF���TL� ����%��ȃ����$���P7���ƖQ� �w%g_��y�݊~�*1�Pͻ���cf?I�~�U�z�"��|����Ƽ�G��~�����TOݬ�v�n�x�:"`���U�wR ��	�?��	�	���T0�� ��u�z���� �۞@ˏ��f�c�n��F���B�L�Fd�x��Wab��WO����L���G�u�g��>�Ir�[�,Q-!��I�6��BC�ݨJ������)���=Ꝣ:���X9��*Y���>��*�ʬ����X����e`��Ʒ���D_�ԟ�����,��� �~�����q�m)$<�&��~0�S�L�x�P��GKv�N�s���%F�}¼o ����pdy>W��!�k�?�ɰ�������~�-D��ӈ���t(]�+0pw`�zy;�d�{��������7��=�z�7��#��ʾ�O������ҕg(k�P��j�$`n��I�>�����{�;)W� �(�c5da;1���a��e-�,Lf�OC+	��no|J܁D�
1�+dF[�;]+���\G�HFsu���^G��&���-�&�z�rdh�=p�]���j�0�U��[�����k ��8�b�;�<��n�s��gٿ����������<M"��%��N6��?��v?v<�Xu�#ܡ��]���{��L>� �5}�T�pʵ�<����7��0z�)��l6�e��'���M,,>��i�$@Y.O ?~D��^� c{�K�ݛ����S7�7�/����K3�;�M�����Ht���'t�����aK/]�c�)r�����"�IfڱIC~s��ݠ�K�r����?�$�xR�5kOY�h�^�A�*����G������;ʭN�7*un9y��� ���$m���iQX� �������G��цS��Z
WA��������3�&~S%���6��O��� T�i{��>��I`Kk*��^�3C�B�lc�O�TE�=�ۤN�hGP��φ-꽓z�]�P�b���O#�3a~�Ԭ��8f�5K�j��2�\60��M�)(�;�D�5r �7� t�p'�0R�O��l=��x�n�;E'�'���'���������9` �Ϻ�1��L��j��֡P���'l��%h��$���I��Nk��~�Ӭ�͹� _&�=%g��!Z��n����4z�>C,.M��X#׳����D}Y1���<X|�"��6J-K�vA6Sy�Y(�����v��eo���HA躚��e)G(�L�.����LY�|zQ�;�v~=�=_��؜�ۡ@^;N�n���?�Q�����c}�X��J����r����_�O��g��3~&��HA��,b(˸�R��В�e<_��fzhz�GA�t˥�cCZ�G� U��iM���a`g�<sGr��0!~<��߀��M<C�=�����S��������0y��>�8��M���P����X�c\ ��y��D��,Ja�_vھ�n�j��1�fQ�_�o�$L��Xj�b�3Ѷz��^W_����Ir�&�t����O@�.	���x�c��̮�h�U�zr�<є�����}W��J�{��" W��$2�,�ҿ��)�H�����Ν��i��q��PP��pHmc~�CV�Cwn@K�#����ћҩ��B��N��t${��������ˮ���c|D�E�� ����4�x]�	������UӪ�d�~M����Yea���Y���"����ߪ����1��60�����(=5�=mN`6��$m!���ϭ��1N�9B�V2V죗��z�9��g
��ǧ�3�hl��ƴ☕�}�;L��#��xXiq�W�0��R�F?c)V�A=<R�C�2�v
;)����5MA`h�>�O��5��[������^�=>�X20jN�o[�R:��.����%l'zy��&���6|Ì�o}����@�} $���Qko��e����j�Nʯ�5M�*�
#���~"�<zk��݌	,����L���5K��<U0�2`t;M���Ҳ~�D 9��nD�o�g���t]���j1XKu
���N�/ݛ.����`;��ǖ�0o�c�_��o���L5Nl�d�L�\ !���!0�$i�NćY��?���Ȼ`-�a��%��t|�.����Q�x�O��m��>�a&���U��Y�40@���7�(��?��^G��m71[!乩�k'h���׮0H������%�`��rm3s��Sכ�W�p([t�	�ƵU�<�����TMm�=>�⹻�N�� ��|��6�.~И��Q�G����u�R:�~���=^�hX�U���R0U�p=�EK�_aX��|�A �yt��:p�|�Q�T�����@Gf{����<�:�q�և�b����[�2�CﳻR��FK�H_D��� �6�k�����k��Km$ v��R�I(ąϋNh6�ʱ3���_�9+��zxG%��/8�~|eS�<���*�  H�u(��!ˁF��b ]z2`�H�ȱ��81����3�-��=�;��9:�ߗ�$rt����۵�Q��q�˫&U �hU���)��+�PY�92�Ѫ\�{I�߅wH
��Ī=���% }�[w��}�*S����$V�8��
N�vu�m�C��9<�մ�TY97@�4�P���ּ�K/6�ּ��۴��(�Ċ��a��P�qV��E.'
�4�ږ�?�@%�{
l���	��k�rZ��D��9=��"@��+���W@��p ���)��߹�z@~/�tD��)�03��N��t��?���_���E���U�~��K�v��6���m�>p���;�Ѷ��[��H�'�2C��+n�⟔~5͢��p�/�u�������!�
��k������\I��8��y�I�!���Y�����/�W���`��%NW�`v����{��*�C~� U�ǚU�����wA��/��� i�j������5�����֯%9�*�&�|�S�a����΀�=M���w�A�~M��7i&�$�b3"�`{�����c`~�=���/D�~����
�X�R$��ơH���8�c=�Q�?��H���U53fOf"7o �4������f�U�4��YJ)��E�Ԏ�ݯ@�o>>5+����U<�:��������W���I·�������ം�w���8N;{6w@6(x�x���c=� e~DɈ#��X�73�k׏� �0�Hj�<�u��U�JG�9?�����{�;0�(5W�х�Ч%)��-�ߵ |5ͫ���'��O��q�Ӌ��>�?�1��l@�Ƽ �.� ���&�Љ���e%_μ���BfH������.��4��%�V	��J�)�w5g�,�4�T;d������O4 gMQ�.���Ȍ�N��5�<f�����{ó��>s�>�:n�Á�/Ȁ
c�T[�{Z�-�	 ��21R7�R�c�,+{�7z�3`h�.���h@�g&��o�7�4Ne:���RzMm*�E@d�C
�����i{~\�U����aa�2@�J�l�� �/Y?Ji���b�2X
6� я��/�(�M43:I���4m@�
��~8G��w��K�=;���Ӻ5�q��)����` P���7ˆ���[��F<��0u�w�P	���
�;'�V�L⦡��s��5V�&ǆ&�9��(@3�<궉qD���|A9�+�V�ɕ�w��Z��I=�����B9���ə_6R��\r�[gzU)3\�hz�����jg�Y���R޶ʁ��AE�A��;\]���x�n ��G|l�(V_fQt@V�z�ޢ	T�ez���_��l_�O�p�!�7���MB�6|=�S?&��R�q9�{�r��u�p�8����EL��h�+U�V�l��|� zRly��c�7\2��`��8U�/�����cϟ �/�=_��&!t����>Ia���V]rf�=X����b�s�l[�|�x��a!��^���p���N5P�?;O��ָ�����*?�iy-C3<CG"}g')m�����wQ����]\<��u��� �0�J�ϋ��I�lWR��º!mb踩sT�|>�LvW#�jB|��w߀9'��'�;�$_t����#j������DT��':���P����M��j�N�J�̂/�b��O���R��kP���?"$����ׄt�|w��{�쪵��I�h���v���_��v�#�5����o�-�oH��{NH�B�Z �()Z�d�(q��V��Fy2XU1_�3HOwO�
�҆q|��#Lމ�ta!q_��$3�T�N��}=���t��	psǄ��= P�Z1�7D ����n8�����G�;��K<`��}.����ӓ)�(���թ�~�I+�L��	�݌���/vE�~�AOF;�pEGBX�:����F�� �dO�=�>@����ٮq��.8�@Kj�3�B� s�mN�����I��RD)1�����0�FB�>�4	1���!�P�I���?�8�A*;��i��|ı٤�b��R_������L��e�iHc���rѸM?�g��H��*��r$���_a�l0�W�B�����8�丫$�����oY��Ot��`<�G��H&���p]�
��o���w�X?�g��R1D�D�Tdg�@=�,�9�p���k䬯~��������}�Х�B��죥�(��t�:ŭ�C��E��VM˻�:x:?j�X�&�;v�`��B_x�sa\���?����s)����G�(*��������s�.+������#4�œo��3��O�����CX<x�d��M�&�M��DmWHu,�a���M OG�앒$�d�u�\�,b6c�&�H;��#S?�Ep�v�c>{e�G��?�s�E8'�F�Oh���X�d�ѬbC2����#����>�j)��}e'�����"��n#IX���9"5�&��l��i���Op�R�0&6 {=8���؈�¨gDd�g�H���O�w��z�uhK4���?�u�T.g+�3ƃ�ƻY�g�eb��~{�N���"&s���p2B�	(��
~� ��~�����-���1��˒��������V*m�]2��C�7�Ρ4���ٵEZ�a���U���O�S�o��n�^_���96c�>��� 0'}�,�slW�U�4|�<K���޽��M?>��`�����©)R�EL %�L}�1�<@�j�0A<Q�Uڇd
����3�� ����LfJJ�X�;T�ނaw��w	w9�k_�w���q"�10څ;�ΔGx߷����]�����<=��)�M�������8x�j�I�Q���;_��~�CY]4HYP#8�k�EV�꺡�߼M��~c��k��{�<y Q����\���"z�t1�:�u�)�y��w����JA:�=	���f��>��f�?�8�5�o&��ږOR���tS}25����o!�M{�/F���R��޻6D����	�f�u_a3��˩H���� LʊR��w����R*~�ԝ\��yFi����A�Vp$���x�uD�"ߤ� �:�pPTuc���P���A#?ׅvQ\^�0�)%�-���(% �.Y'��\����`B|�l��㐱sz 1��_�OD�ǹ`X�/IG4Ғ�j �R�ɫ���j����&Omj��q-�<�XY�:!th5�T��O9FZ;���h_9�s��<������'���/��E�R�O7�.,u痘J��a��m 6u_"�pVuZOήѸ�E��sK����ބ�R<�5�7ࡃv��')xG|�,%��?F�h7����|�0!hQ��b��R��j�8�U���ߧ��m��{��1��g�+�$��{\3k�c 畫P\���""~g=�W���R{��Ud�����k������M��T����lB:��;?#�,��z�O&����Yfa}�\,k�D���*�m���FL[�(����5�l*��SLF:^���D��%����40�t�G����$�Wy��V���G�)9f�-!EGd��Y/'B��/WC���I��N!Q�|�}��������0��e�0�5ea���%*���Mi���J�tY����`��['��lF�|� `���(Ǆ�}�4 �:��ж�i7��=Q�������R��wv1ט���H�|�ҁ?͈�e/��mX�9�ڦ�x9�{��K@&�,�,��'��m�KO��4��5{ �(�',��˩�|j6\lVk�a�?,�;;G�P�S��/_ ��0qE*�b��Akx��g}���*���
Ӛ=p1~�g�@Y�z�]8\�6�i�/��Ã!fp��X��nώ� �i��!(��������Ys�4�iĿ%�/�z��g�t�[wb�I��?1R�k�d��Ab
�E�I'�D��ͅA��.d� ۲�C���O`�߶L���������r���F)	)=dh�F����d7o�r�Yʹw��aA���i�\H�QU�����%�������;��+5���^��g�
��7��K��ހ����()_X�K�#Xdoj��}]1
��YXy��2ā���(8��+�f#�NF�9K3!kg�
���oA-��`�����}�A��	��F�st��*��p�����:/x5ł�M�)%t�PJGO{?��9W�*p]L�юԘ[�����O��o��YV�젃@1�\J�U��,�dԒgTf��tJ?�悼����U!u��m�٧��������.��Y��T�C�B���G�f��v33���F�?5tHԓ��7�S��P�"��Np�rG35�`�&i-N�w~���y��J�BK��m�u��N/l�"6cE>^�1Ȃ�����X>�)HVA�G��e��:���,�75�&`����!��S��sr� l��x:|ʫJ����WD�V��$@�O��d��W�v?;o��Eڶ����2Ƽ
7h�#� #�c��"��� ��AJ���mX���K����ѥ�Q!팋pA�۵�%%Ԕ��RVH���=ղ�-�|�N�S-�-�+xx�H9���3{����س
;v�H��<tl��!��'�,.էFS v/�'�#��p;�n4�j������X�����%���|U-�� �����).+>���8�����t�>"��x���@�,���`�F 쌲�Ne�%���;�d�ibA_�/�0���O����oQO\((���v	��#���X�`��L��������e����;� LQe$6�Y>XO�ݯiD�As��xQ�aő�e���ؓ���M�A�wQmvz����*�#�iRԕ�Y'�G��M��F���o��Xmz:g�*�T���H��ֺ��wdE�.�X�v(����Y�ȼQS�]u�0qA�MCz���V�o	2��:k�p����M��F<E��@<�<O���,l���?�ԕ�иY� �V�#�ŭ[�Pl����`ZZ�,O\r��˕8MV��ޮ��6ёB�oRi98���9�}�{yO?�Sm^����@��W�����y���M��9�̖�V�0>iIN��Bv��'��Q���z�P�����
5z�"�?�}@9�u�s��d+�X�s�7Y�O,ĊϻłU��Z��SV)��#�vc�`!��.�*�`z#~�,k�~N	'%1�y�y�tJ\tV_��qZ����q:��ld`<����ǱJ�kSE���ɵa�a��wˏ/p��q�� G�=�?��p��!��-I����>��h��Of�Z��l��ܜxr��>�y�^��g\��1[�W��c��i�m�wP8L���׆ƹt��)�H�>  �������SL�Wk��E�=��H��L �%���Ը]��»�d��|-~���C0M�B������\>�S:�(������v��y�Q3A;��)�����$���ƀe>u5�<@�֔F�
`���|Cs�Ҕ��j�%�Q��c��e�'='�2k��+��1���e���:���1�"�� ���k�������dS��Z�f�n�y5�� fo�چ�ln�_���]��>�z^۫H1G�z�z��9L D1��2W�U���Q�|��]��(;�x����Cx|���1����SG(`�}�za���f�"V���E)��W�p[O����hr��jR&���H��)�Wjj�]�����G!äo{�;~+���
�B�N�@	f@�_uv}=�L*AJf��_aw��]E�0��������ļ�C:��+�P�SS2��>a�T0|�;Й)�s���de𛬔�>r���H�Ɨ��+C�d���`	@�ڝ�s�Ưt9'\6�ę�a>+��C$���wHo�����'�s@�M,���vV�����
f�����O����@|�U@QN�މZljh�n�+l�*�S��Nrjl�0���F� �ȝ
��No&��� Ǥ*����lV�m��a ��K��́Oy����޹[~���-��x����<lFD4��q��B���틣�G9
�Y�q)6V����}AB�Ч�28�l ��͹8
�74I����
V_}������P𪞫�2�7/�g@��ԏ�^��4*6���V��L��qp�R�'�J���TI�=��5wf~oon�i��������ne������7�T�g�-�(E�)��Ww�-�M,1�q�߷ӽD�U��m-�ҏ�ҏ�����|`:�HW�qrdU�P� �ff������H�]����F��n��x���a��]�"��5�-H�|����܃�J��27�)��9��We�EH��S�d 
���S�)hp�������O����s���S��h��p��f.Jcl���7�|0�"n��&��dM�O�=^��#Pp���66�lL��_�\�f8�$l&-o6+
%9E�x�!q�Y��,�ۓ�{�lD���r��ltw��Hw��.�	����?j�Ǚе�+�}\XH���i�C�t�!�B+tZ��?�0���T(����J�#;?�&����\e�����AFj�D���=��)H,�-
j���UR~e��t�6�J����8|<�tFo�]3Ézt9�;P���{`��XQ�WvR����!�
0���>w
<RR�P�ֵ
Dod¿�#>T6���q��c]���(������ͦ�g�ݎ��e]�ŚfO��XLz�ErES	��f"�#�~�����'@��3���:��%�/$�@yaU��[���;��w�����]bz��<�X�<����n'�k��%�Gv��G�T��ЛE��{w~>��$�@Z�.�0rE]��U�<����ݡ;�YD�|K�Y�ݦ�:ֽ2o� �"-��]�E�@k����Dn��"_}�^"ʶ2����J0Yg:���Յ�m��r�{|7qP�#v����ʗ�?�{����~Tp��b�b��RW�����.F�m},"��:����b���
N~�P��
m5 da��M/x�[wn1˦���G&�*hT a���5 ���4��'|��.ܬ~<���Us�eR!�Gc�Dur��%N[1ɀ�����W�e��u�b���{�#&���rƏ��#D ��� ��EQA���Ua�z�������1�4�l�۩��v��&��#Ne檭Pej�]��@��`��"�*��9*�0��w:K+����@TD�U�����y�p#�G�#���ĉ������$(bÍ����ThSMmB_�UO�9Wu��f�:�MN_My���G揑S��F3�Ǐ�����Ϲ;��i�ɠAf�Rk�9�kP��N&�L�����x�R�åF��vd��}ڹ+����?��x^��؏�ӡ��ް:"�:+1e=,�;��^����@�V��� 4��;����?�E(n��7�����k7	��:�ؠ+)w�^�b+��cT��
>T��9�Q���Ѧ�._A�'?�iQf�ی���p���>����2��G B�0�Q����#��#j�o�����4ړ
P��R�����B�4k=��]Zq�2��h�OP��(x �'~�%ޅ58�:��Mػ�����P�i1
'
i��*?�m�yc�V��p�e�f@~�\��e�/-��@l,����&4z%go�A�:���>\&<!"���P�� jmj�����Q�ȫ�~(�`װ�k�{@�Na`��Qߑ�:��J�%�z��  �G�Dk
"�m���ԇ{���v_p��5��1��d��4�d�@Y���M���m�ǩ	zc���$9P#�Cƴ$����Y�T�t����7�/@��'W�Λ�S`G�tK��.')ˋ<��'So�X�%.�NȀx��jǂ���H��F%���w.J|;�C�
��)n���s ���%K�aXA{6�aLB����i����b(3E�yz�)i�%�Pd��"��0����o5��)�]��P���hLɤ�]�@m�wye�b�hM
��F���V���9] E؄ ����u[J@7�lĴ'�a��z�s��;�7�%d�>��ϛ��$I��D�X\�8*)H	�1|i>J$_T�ٶ���fM�)��L�g�(BW����IB� �*�
��y\��  �7"7�lH���
��@�l(%�ڭW���`��	�ڟ��Ek��d�>ɯ4l[\���������j��f���^����ŁT�[MB5n���H&���:%��Л��G�L4��p�IU�����id��U�b�u� ����$e/�����7o���r���*+@�|��B.~.�c�8�9�F�$�Tf`8��MB��w�P�br]GY�H�g�Uk�_^�����^�(�C�ĥi��kFnYy�����_y8&��w���W��ع��<��F������xM��Oz���?�86�R�_'>���������2�/)!O
�	�'j<#��ۮ������<b1xY�S��*�fǝ0�+�R%���_U}�:A/�K|JC�ˉ8�mm̀��m&k�`����wadÖ��#N]c�~��y7�4�u��턃�EZ��J�̀qQ�.�@<�SF�˦;�h��S	(��dyo,�ྗZ	��9��4�A%g���i߸��j=�uD��`3��@"?c��}��vu�<J��Ԭ;ѷ]Z�>��i�s�C�^U��|�/�k���'�aߖ���R�t���R��ovo�/^m+��f�u��ja�Ɉ�wA���"(���\���'�~dŷ.��<�6䳿C�����$U�p�e>�w?'�=�V�����Ɇ��Z(}͋[�M���B^��R�x���ë���,������k)5��n�L���.>4q�.�G���b�����¤W��4ͯTҪ����5�I/K�����5e�w;��v��>+vI���E���UpPu�K0H�e~+��T�jGBG�����X{���	z��3	�؛B�0��AI� ZR�Sr���+B5���<)�ϸ�0�dTRN��5��捎�x9�n���W����f�4���k�f��=3EPFkU_�g��m�]�u�*7�I��S�t����GE�/�z�d�ob���3����%S��LS(D<7�"<VK1H|�׎�6�_�9`��uNk)g��><�@�X��ߔ�sE�_���Ӱp&�u�لZAd\�${�M�����i�#7����J�Z�g�= ��u�"<�[��������F�:������iȼ�͉Q�V������w�}t�4���z?�N��t����.}=}��f����>�F�7q���U���-��Y�멲��Ǖ���*�ǎ�Mk�+-ʡ��=��d������}�~j ZRj�;����;u����X(|�K��!Q�1��0-�L�{gBTH�b}８�\�����'�k��7�;�G�hT5w�Q������H��t����P]�h��P�n�/0o�뇭c�(l��;����o+��lV�V� ���>���n�qBxL_�Ff�ɉ4 �KFr�Lj'8O�W��]�՞���hK�y\E�.n"��2���m��^�����������D3<����rd1�|��_�c�<˫-v�UP�*�B��o��=�{%�����~�P��V�/�}�$F���;�<E�_�=Y#��������nm"�S������_�\����b����E�{��l���s�I��\Kr�`�2�uq*����ڂ Hk����u�	6�ڂ�ػ9��*���S�*x���9��R֮��xM��{I\��M�w���)��斪�磶l+Knq���"��XK���#�Sb>���6=�ɱ��B���u]�P��7m�Az2cb<���߷�H�Zy��SJRR�"��/���N/��4�>9C��5�˺@5��[�w_��l���仅������|o7�3(Ȣ�c['D��jb�e\0��ɯ<,�-2Ɗ��w������g�j�i�M����3{=���>ҡ�&z��Kv�h�F�҂<]kY$�UF�:|p�B<m��106�:e�z�����(�0�6�L7�F��n���S�{NL����X͑:�s���F�9�
u�|Пۙc��G�S�M=�>%8��Ļ��i�#��v�A��pV���r٢��ӄCڬ�٭l��b=��R��_Fճ�zvϢ�g��z��.�i�g�������Bh�m��{�G�D���%P$��8L���
w�S��g�˒F��{/�̙�]<h��ر��f�&�]5�oC�|�	ȥs9��VT�������q���������G|�z�m��8�������/r�ȝ]lZ��
�珉�'�~n�?�U��`ɕP�6��G3"A�T�/�~�1�V�`&�[�~�r>�
@����xD�v&�`��0�ąO��E\N�'�`gc�[�:$���F[Gwx�C3ԕkl�R��C���>z��������>�Վ�M�K���h#����2� �u���`�o���7�t�ʳ.��{�h�;��S��+I��Ѓ��e�����ܐ�g-Ȯ���B�},E��9.˸Re\�и��R��˼��T�}|�t���ӱ����㗙x(���
�U�p�(h��c\s���c�04K�:����<����Ւ�(~�7�=�>�r�B��[?ەB^\���?f-Էu�o��IP3�s�yU�.������[?gLt6�3$�������G�@7���<�f3��5���[~����z��	��J:�tU㇂�����Źz��Z���0�Cm�h�O	:RM/��2���_�A\>7լ��1I����g�u�>{˓��Ia�Ǥ��'eo>m�o]�)��y��br[k0J�?�g�\�A�8��][i�AJ�J��=ڟ�䆔�[3��8�C Ay��"��bF�(=G9����(>��;n݉��#��H3v��K���B9�P�N�;����d/o:j�Rw�xSYhĢ2���tl�nHcUX���݉���K�t'�Z����P:�2�w׈~�:^��8�/��&XE��Yc�-{���i��\ѣ���xS�g�$��͹��Y�4b#«�D�ݒ���J��5��٦���6I�����ȉ �N�������t�C��z4��w*ċq�#y=�ǜ�z/n{N� *��]��F�-YT�^�ˌ�qS���{�/�9ʋ�=�D�O^��V{��b(�PP[)^[����)����	(PE��H�`�v%T3��/N���o���	,�*����Ȓ���>zъ=1�J�\Y��e'30S��?��dƎ,~�" Z<t)�k^y�i�
0Wإ7�k��)����r����Sc�pl�WLs�.��j3��.?];ѽ<�Xle L_ݪ��4ȻSf#5B>/�&���X�I�]�R�a�ʜ�C����P��w�f@�^�?��BlY~�'���\�h��]��"��6���ʤ9|ns�Q��D��De�;�a����ؕe?����(�?��"rĆȜ�T�֭��m�sCIo�Ȫx;:�'��R�X���3"Wƚ�N�\I��UV)��kR��<� ����j���:���v:���S�L�������W��w��^�Ո��O{�/mM8-o����O\�	Q1$�Ë��шTqb�:�ٍ�N�8�Qac/{4���w��d-�A�2�h۝��UxT���2��N��}�+��Z���ZPM���%��j��$ҋ!�n���~;��%�Lak<K�򪓨%�ޝ�*n�b
�L�����NT��ȍ9�a���\��:&�l],a}qW����?�;ڷ	�����H'4�u�y�wt��/��Il�W&7�#�s�x��U��	���	�un �a/[��#]tJ�/��G#����!0�}k2�S��ͯzY	�&U�.X�Iuh!�i�+U��Z~��#��,�p�T5;y\i��|�<�}@N{|�
]�r?g��B=�r潌��!��P���鎭2��s;$'&�t[<Sa�U]�+R��cZ�-���6�h�8X	Ce���	����d���Sǉ/j�u�i-��s��tO�kH�i�Be�ߑ������,���;���ߧ`��5�iӖ좹�����pn����PHV�ҟ���!��S�RŔ)6pۅ��h���b�	�p��#"W��#!�d��\[��k�������	zz89����_/��,g�N�=.��R��R�¢�֏6�1���K�����С$k[j��N1���F�C����O�)�tJ&@�!�¡_+Q�&���j���f��f�<������:R�>�~a�P��o���T�Z�,��pwe=RoHW�U�Ђ�T����C�g���%&޻�o�$u�ds��Ea�)��4�0�.u��9ؗϖU�����1���W���gs$��X{�Wڇ'�+�>��y��W��-S�:�׵j�7���!�:_N�*�Z������YH�2���|4��r}O�i!���1�q�>E�^��c�hq�wڌ@������R�'���3ə	��p� ����ԉXa����7��b�vɓ�e�X����O�L坬�������f�!��H#8\�ULMTG�+�C!o�1-3�F-��H`�M�h��#y����4G����^E��2����e���G�50Nع��7�c�΢ӕ�\����M_�=�����N���7�c�D�m�+$��,(6�6�[z��w$���l���$J�7�{�+��q91��^�iV��k���ap?J{^���4�%g���Da"�;jͨ`dH���؁�G���G\��4٣Ȓ��Q�G�-/j�tf�%}��Ǧ>���x��O1{;ߙi�
��_/�C����ug�T���a�{�/�P�����������)]�2W��������C��%20L��bb/�/�2�p w�娿�3�e�*�R ,p8]HCۚa�l�xw�$b��!��=`�������1�o$A�D���*���IȚ����Z=t+˦�"���䗆�!�%-&��XѦ�agQ��}��Q���> <��� ��G-`se��l�B��օp�e@6T����h�Å ����2�[��2r#�#
�,mp�Z�t�O Aqe�"��c�s2&��>�[�������\�z���	��R��}�6��3��XN~�>޶��]oz.��p"�J�����V�n<�L��v�����Pk�V/�����Ҏ�z�E:�4�erC�8-�OJ�b��2x�/z�
Ͱ�Ŷ���g~�0�4�<I�;q�{2V�Dj�a�i_7	Q߾���b���ʲFޜ��\�F��R+j�@ A��W�)KM�<i���޵�d���duJ��V�̋�������<��m���s��\e�\R�tl�����QRR��k ?�r$Vyl�@e�:dd!���Oh?ͩI�g�8�s#�Er�A�&��S���+{S���8>�
9Q��1��+Z���x��������t��Q0�i!�����V��d�z�涴Ė��:��V�s/<��N����A?k}���:Y�y�zפyӯJ�9���'���Ӿ�K�nǑJQ��T����x�iQ�������*�	���Y�'����kC���Ƿo�T'ၶ���p�����!9��K�l�_�٫!�"����Ԥ`����&@/T��exq��oȭ�N=Hl� -S6���0�J٥�)[���%=�������8����S��+SLV�!��)��%!�VQ�!��6��5��sE#ǵ}��:ޙ���k������KJ8�v�3�v�
��׌��٫��lj�g�������-?+�[����J���˻�$~-�%��-���_����N�4��j�^�7����㾩�PEv/��+���O#�B?��v�4�17I��8G���D�mex�n"�4����[��������%�(��Z\�,����^�r}�&Mn��6>澯�8CO��:�
�n`��!�V�-*��|�0=�����y�s�?q�{���R���_��k�0T#ޅq�ƥ�|�$7�r,��`���_�sF�`T!��Ý��]ա�`Eٴn��a�u�1ػ;]����(����､-���z����|����R�X���7΄�lbyŏ��7��~e�s�D����H�p`�l_2�y��O�sݹs(l(@�h�v��a�%as>��3	v�f<�\oqA�ށW)oR|y�x���w�1�ьpcs!=5��G��4��
}����t�RN���Ҟ��s�����AZ�šV�%����I-Ӯ|�D�tl���ȭ�W�V�����"�G���T��w�����z�A���5�ʁ�h��TΟ
u<@ma<l\t���wO1����]X�󩋝꟩��i�8�!R�������?�2,��{{ i�n)A�n	E��:FDR���p���!d��;�3���_�_$�^{�uǚ�9���������.�鲹~:���ʪ�����/��ɠS�y8��R�g�%4�VN��5}��\`�S{3�(�8W����E���v�*9���E.V��;dv���)^g0j��R��:aG%����A�P���P�^��� �+?�+�e� ~�:g�� ���N�Q�;,d^���PvE�bW �]Q]����>P�n�E�I4�}����h�<���%�w���N���K�%|�"����pbW*�zB��@�u��ɐ}[j$���o�U彅����uSCtV���37�f���z�
rn<���g1�ȴj�=����D?C88�{\�G��ۀ:}'��>�s,�䁎Y��] )e�Y�V~7"���e���Ϫ	��L����^��p��-�HCh���u(s�	q��s������c���Z[v��.�]���w��P[��k��I[b]X���L�+A`�,s�{E�`˙�쩰`�9�w2�q��[2:�B�#�r�q?�6}^�^v�.E������oK���g����a�{�fJS��
�������=��|<?�-x�VAs����ճ�vGu�8&�2� 2vF2��U�@��;���X����|�J�ħK�z�����y5��3^���l��H�!),�h�E����1S�dH��.t]F�+ey�(ſ
r �6�9Lr�����Lt����s�I��;ě�h=o2ء�}�vW�_�3��~�������:*�x�J�.��?�O$�L�YM��.�;��\	���1�;/�9���i¢�k����	#ƊV47��D��/_���[l�n�AFs�x};ᬇ>����S��4�]X��i�u�|ѽC^^�kG��3r�/8T����=�Jγ��@2���3�D�A]�c�!˺�+zkB�ì�*|w����)R�M�*,��fO�+��V���&�+@+ˍ�
[xH� ��^��<�֞B
-��dU�[��w����ſrpV�����w�q�i�W�SF��~3^�H�l��QR�G�+d,����߿�8��/,�_B(ܮt�����7j��Z��a������{�M��.V�ُ�OS��%�V�*��+�g'!X��jk�>4�绂o)�،~q���H�AZ�aL�5�Jxf\�ט�t�	�J݀^|ы9�GP����ge�ɬ�<�8�yQN}1.)���OD�hd�Z�p�Ob�W�22̕(��,��P�ײ1-����|��:�A��t���1�paC�7�e�@�2�k�(	�W!�2f��ڰSY=�$��~f���-7��ظ�h�p���yq���%���H�E��j
ǒ$נ�Ǭ��$*z�y6H���_���M�їlu�Dm���p�IvZ�M���0�"D4	�K�xɈ������i�X����L]8�}��Ҋ��WOp蒅��0�R���ߔe�vp Z���^X͉�y{ǊDa\Pҷ�5�<��G�9��~O�A�
� �蔐fh�u�-`�Ȏ�ʹ�c�n-�۩&(��,����Q��C�ć�:G7=�k%#��<�W���Y[a��ơ
۶�vc Y}��[��[~�\W�m��Y���4W�}=�s��A�ar�'�G�|��DA��tө��2W葤�}Or��s�r�j�r��k�����0����>��r�v��:KYg�����L��uA"��=�3��F|���.Mi7,�t�tɫjm�N�f�b���qM]����#�Gr2z3�_�,Q�a�f��s��@Gn>���$7��:F@�܍�����l�o���N��|��a���'��ә���Yl���2sZoF�[t��P��Ք�<�c��
e��G|�x�/9`�n��P�a�70��5Z�Q'<wΏ�ns0����ĝ��>ƺy��M��涪~EH���+Ţ��Δ(��ֺ؂I�brLc�oq �\�Q|%��Ʈ�u������j���t�����MWֺ�p�����pCv�r�W�_�6�
�f�-�_`�����"^�z�������R�
o77-�B����[$*Z��';�0�'�%�9����ہS�l��jn���-]x_d���1w�V�]���������(�O���'�v����TH�{\T�9&�J��Ɲ񴼦�¿�/�0��_�ا�;^��C��.V���$w�_����t���`�~?�c�S9P�Ypì����cD���i\rEjZ�x+%�0g^�n۝]�Rfj`��FA�HW{2`c��i���A�A�vU�V�v?J�AZ�g���!(ԯ�y�p�D���MIi�p���}zu�W�ޒ	Ɩm��^��b6؈�GF������X�#����<��蛍݌�C_���u��G�,��~����ma�LjOr���t �=Ix�Z�� yM�p�KN��1 e^ګ�|�,1�g�dK�����z��6��_��Ҟ<��_H�G�V�����C\�������f*�?܍��b�0����/�(�\s�5�O��8pu�ՄF-���M_�J�h*�跟:�Lz��#�C��T��2���,�ء�UB|��5�_-���%���T�L��ڴ�|O��k�]c��ɑ��'&ny�EW�?m�H!O����:7��x�=0�:�������UI sN�3�M��,��oq%ԙ�W��h�T����G�E�-�Z�j�X��G���P"��~0+
��hP_����x��@=�+���������z�噆���<���؆p�����$+�����["�|�
1\�l��1*%dl4J4,�6#62��O�7f8]z�8 �#�	� �����G4ԏA�5������+D�Č^光�'���z�h������'z]hU��b���i��9c(ܭ�Ok�p�7�1�/B�8+�S�=�dK��X��+�J�⛘]�i|��IZuX>���2~��zi�^直S����ʽ����B60�#'ϣ5$�Ҡ��1���_N��E>��hY3��R�g��^��G�`K��ތ��
Q6	�!��?�ң��ٶpQ�vp�����B���Nګ���})͈�l�{��N�atp�۲"�K��}̶HY\){��C�MT��ηK�
�W�����*�
"A?�[��l{��F���Y����ؚ�%uf��݇xn���S"Y'z?l����jy Zm5����2#��P�ˊ������{HS 2�O�L�j2�"?�Y���œ�цd�@A[#*�स�6pb�����\�ֺ�,��)����j[���o��`tO�y=�q�{7�t�Y���=U=mq�����GTJ@�S�jڸ�����#��%��2 �N��������P�F%�}}�	���FQ&�����lC_Edc1)��B���^To;��K{ `6�b;6e�������Z�(w���x\���w;�`t��I�f�ala��`/p�l&>>-�����orD�����?��2r����<�Л�?:���uC1B�_Q�B�2��Ľ'�������RP��T��6
�Lb�Y"��%��m�sAX>Y4'� �>��H 	/�>	P����j���VWM���4������Ι�x�<�%�]��L=�
PB����pw��I�;:����'Э�v§G�&��W��$���"~�SVt�`�+{�%O���G����'&�eT��b��JoI(W\�ۇ�i�!�k��'lG?���W_[�Y8�}sR����X�o.�������b��*���/a_p&y�7i���~S�$�5��W���>{��S�`BI�'.D~~El�͂�j4Q�ǐy N{��T�Z��@�&����ݘ�M9����,ӡ!�)h���8L�&!Wǐ��eC߾�L����q�燖A��[�,�{2S���!_+�L��`��b�x�\�|Sv9s��N����l��2As
WW�	?J:b2]��<%{�ǰ&�����\ٿ��}�;3�l~���!r��GC�Ȼ[�W;8�����LaUb�Pi;a~�L���|l�r��Y`���lٍ3�w` �ŋ�\��r��N2���@ά
v\,F�OL+��li�R���*ʸ~a��
$�`f�Rq'����6=��g�Zy�qOwj�D�ſ���r��E�,�{;j��g7����k1o�6�T��P��y��O$&�����Ipo��2��ox�ZҀ*�Vӟ ����M���J�A����&3,u'	�� =���4��]�Dx g�}�.�[���͋�Z;���"":S�J��0{N,~��Һ�B�g�sd��'��UL%8���~��E���r���81��� Ij�<�����.�1�!���B���U0�r����r6k�3��֢*��O�d������l�Q2�v�ˉ�P�D���B4��n#ꑜ�QK#�Y�RH�/���x�b1u´�w���^�:jB(o�W3g�#20ɕ6�R�Ÿȩ��^�cЗ�o�c�,�|������5�l��{'�@�#�cd�Q����f�oVS:o��"�}/��PE6G��X��m��{k�FXEP��e�qSR�/�+��v0א��M��x��ߦ"��S�k��AԄ�$a��u/f�b;�2�vw�v��X����G+ݍ���Ɓ:-5HN��]�x� �TU6�Q#�H����e9�5ӷ:g�HB�e��f���F��Ԙ<��.bvE��z0�	U��>ge�����*����{@�ף��~��ss�c���EP���,�X�\ɳ__���+���@%��_��]���p�?���U@F�K��k�G"���kN�f�K�I����l���m�&#���q`,�_.����>Q�	/����A�*��/�m���Q�o��/,�W#=���0�Ob8�eX�k��iW�R�"n����$�i��Np��F�?>�`��6���(0�b��c����#k�0i�E�X���j�^�;D��6�Kc����]IC9����w��r� ���~"�k�V���K-�N
U�	¨�?	Ș,T@`GFiV=	Hc@�c_vM�:�a9!:4>�<-���� gE]�Л.���^ԓ`kf
iS�]j���d��00��&�N�	:L�?*h��(j�5_��	�5 9���n>1�=}�M�B�8�s�!ѫ$�k�[�*%���*���&�� ��c�~ŧ�i1z��]4����N$#+b�`e~�Ú�v]�WK'��ɲ�N�.�͂���G��$<Y�1g
c���V
�ԭ;�H뙙�F�I>˒i��5{���߅	p�L����|S(�����`�.=��
�܈A���Y�\���$Z�۴������ތO��s���A�9=8�~��D)Nbhby����B�w:fA�O=ċ>c��B��������W4ͯ����1�������hg�;8���M�1=�n���.���~�����4;�m���Zm�(����;a��Y��O�X���[Ѱ<�V#J�a�P�J�㮋��JfA��c�}S��g߮u�g����Wi��'�+9�=R���i�x�T��F�ӹ�e��8~fW�ҳT��� -��J����2��O`�M�h�[��α���KO$�hԁ�Jc��0��5�w�������ރ�Ɉ�t���v��	�mU�'����c���{�@����%ѫ�jm���"a�%׍�LDA�,��v�K
 M�U4�Q!�\��¦��e@c�ʸ�o���w��͡������/�y^I��b�s3����`5*|�.𙛴����=7���&���l*�����4���� �$����Ƞ�8p��yU-NF �_�,�@P��١Aƶ���(@"��'v5�C��B�����R+�^��eF�M�o:���Œ
�F�g�=�d"#��1�)^L�@��3���������t�,��l��HŒ��5�B�na�?ї$��ser�G���_�~�k-Y��`�0�QQ?{N���n("���$;|��C���u�B9�;� �
�PW�����S�Oaw18�-͏��]|�����k9*J_�J`�T�b�yo �|�F��{55ܼj��K\�|�{�I��6l���
��bX��P��o"�}OY��Z���q�T
<kR|��Bɩ���!�Y
	��z��9��RW���(��X'uVKys���z?�fH��zy�����,�����e�ël�l6�B�����$�g�C+m�[�k=����(�s�����G������wo�*n���g�;878k��
�g��w���o7L,��	�[fF��N<A!n+�OS֪a��rd8���}�8���~-vzwD!����Wc�6N�'�T�;�W�-����9,Mw�Ӵ��Qb;�N;*l@.+Ș|<��oS����Ŵ��h����=X��,HC��SG"c>����K=*rЩH=������[�Έ��;�4�V<� !�!����:6p4�ԨGx�*ж�]����dH,������s[X%��E�q�D4�i�{s�W5����$B�;Gۘ	&��@�LqB��i�DI�;����ۜW��P�4�8�]�[�b��}x��W�k�Ku���S��:x��/q/e>�1��1utC��E��O+l���~�1BM.7Ud�$� ��4j�w�&���p�lÊ3�R����r9EL�P4hiD1U�X3;垺M.�;:
��`?��c���K�4ش�IQ�, 	�|\K��>A�+@5���3���m�SQ$�"ϯ�fC�
��(/(5�睺r�lT���_!��́�=�_�!+i���W�<��9�6%p��-*��ʍ��F4���W^EU����HU���j��'�B4�lpM�����-�����F��[�(e�[VE��:X��9����h�%T[s!�]���9bB#@�Z[G�9\��cEȷ �\RGKԚ����޺�}*��G/���D���أ��1�w9�����_k����
�7�Y��7kP�B���ȽJ�|�$���]ߋ4uuK8z�~D���92)C�u�޺[p�"���1�+����Ά�$�>8TO.�{e3q*.|�����"{�w�����=	CK�"�)�G-�g�j�9 �R�&nF�T�
ʾʡb�Y��܁�A*��`*ǀi���.�t�u|����q��7��/����&6�� S/��N8��}�f���;�I��=a��"�F0��,اX/��HY���쫆1Gq�OCi�� A0���_�������n��	S�����D\<��t,}m�����𺭾�d:X�=
0	��Ś�6�h�Y@`�tYMC���$�"��i�M���/"}�(C���R���bȺ/�;y_��F�k.��7�v�2�oK�4?��zL�6gS,�4�=w�}$�@R�0]�2����OwGF RN��M2t�v$m*�E��y�k����
O��e�?����q&Be�3nf@�GK0�̈́�iG��`cz��؟ ��/rɭ�a��\���������r��"��A���/y1�>�崅&˂7`U4��M�s�s��u���Zڢ���4������q��޿�Q�:R�����`x�A�����c���䯛w/^yh0�z� ��ehd̋��74��$[�IjX�a���S.�t5�>�~
��	ܵN���1����^����̑�ۨ�&����Hc$�NJ�V`G�51���(*˛WA|7J�����=�G�B� ��Y�ѵ�Q�z��h�+f�r&���}��{v��5�>i�:���&���]���%F��Br�ɺ��Òa��'�'t����fs[F;d�HC��U����Xb茥�)z�!}H����;~E�Nz,Ж ���Z�#�_���pA��/�aO$�"UPm;����S�is�t���Mf����̄�3O~��votĢ�G�M�Z3�𻟾 D� �Ԍ�~�h���7EVw+�P�L��X^�Ѳ�����H��0R����{xP����X	9����pMPrC3��[U��׺9��F'!/{T7"�iam����Ź9>^�ϛ�0T�+oC��?t��s��Ō>�14M~+��'Ҝ*���ƀ1���+DU�․�_7Ph2��$@b���������)PGvJzd���ű"���zG�0N'�;�<ک�-��.t�&q�	I];N�J�{����yi%��tT�z���6�w"�O�N��.�����ֲ.W��� s�?)1N�^� v&��Z�Q�ŔwC�f�g07#ּ�)���ڝ����^��~���o���ħ��u�W��kz���g�����:�zt	s9{�t�-F��&m��N	��[�|9����4|M�EA�h�*�;��
�l�m�-+@6sgR�0��W�\p'9i-����s;z[)�����G���_�/�lun���㲽�bq�N�0��q�XQU��i�n�jgݾ��j����[ �j3�F=���O'���Pb=2��>�[�/�w��%�z�LAH|�9B}&�$�,y��p;,I�u��@1��Y�-�q�O_z�V:*��^c=]U�fLc+�\z��/J ��VϢ/��j��Rnۿʑ���_�7��>Cr����φ���GS��4ɖ�`!Ń�3��6���1X�Ӌ�D��A������W{�to���Yz)ʞ{"8����"ZxLO@�U��LS��Q}�8g���>��`�/�m�Yꪾ�*���k��)����7'6�A����tT��;sHc�J՝��%0�Ⱥ��x��^�S���R\<�̻0���>�G������Nv�ʦ,�;�b�b�}(������P�:�b-s�0�l��豁K��f�n!JCn����_��@�mN;�Yj�}���y^�TLf,CZ����+x�큨��*i�P�~�/�F�)���?�������J~�r�Yd�����>�
RfД��a���mq�s����YlDg�?���%�XI�l $�hcK�����������J"oV�oZ�̊���1��pX	 �C%�;?]��g�l�!4�j2%�^�\=F��U�ثq�QF��(Z�rKS��(�Բs����H����ו���:�/_�o�Q� �6�[����f��y��w�z0*���M# �AI�5"W6n������&GW��rp�f��w�c��~�00*�R�b�xI�>Y�����K�YN�7��zސ��>�2/]�3c��_���w��)��	��>Xg�t8��	1U��}��眨��-7�9$F*A"Y���Uߦ65 c5nB|M�稞hh0�w~۳���#:�H�����Z?�U�uLD.H�"�!y�ۘ�K�r�qy�>�c�?��o�а���_��\�1��& ]j��ڜ��=$4�E�?_��)�J��j|��Oc��k��ꇿ�w/��Y����V�iZSyL����V������A6�OL�ꭓ1�=o�\�uQ/��Vﮊc7Tz��ڒ�
�5��Hi��6�A���Q��X|"g6�sׅ�0�=�P$'��+��|�8�W���~.�I��O���Z���۳��(�g�K"��qL��v�ۻ��dV��4���G������1��Y�2*E����I��3Z�J�������#!���R�l(��6D�k�<��d��\�z� ��'[�Bw�����H�����dCP[3�<�,M�D�ǧ1թ��ʅ�Vy�q[�il5:)&�aL$�J�*PM~�j�l��Է�� 7%�����?Պ	��r�ucܣ���a���U�L/�yF�X���.�y��MA1��K^���$���s��=y�<�!�SNyG��5+`:fr�����	�oU+�-\.�\��z��A�|_B�����r�w��<#ƫǌ��Z��lY��?|�b��.,5�!�7�kU��`ɑbk���0k?cD�m�,3����b���E�^�H�`/^����%Nz?�ߜ��T�m�Q�ܫ"q8�o�b.-�D��n)������0�f�!���}2%�zN���G����h�z,rU�N�b�T�� ��<��8�7y-����Bd�+�9�����˾n��X��i�*��̄�
������3?�!�Kv������J�H���>E�,Ϯ�􅽈�=�I�u�'��:�q6�xl-�):�̷ͪ�Tq�?��6C<u5��1*5ԝ�6�@9�8p�6�hy�����'Q�7¢�l��-6q�N]�Oڅ"B-��z	�Z�s���Ƶ+N�ĩ�ĸK�0��M�j�f@"�*� �޲��2�F��rE�%�U����Py�I���s`�߹��[�� t�����΃�ɧA~䍹�S����2��F ��g��ЖJ�M�s#u��(���������r�`<Tɥ��'k��u{!��e�� �Z�g�{,��m�\G�s��,K�D���Ɛ�߀��{�����G�i$@`^��1�ѷ͚�Y���i� �9}P�@�Q�1��	�a��D�1����e�/��1mRޟ%��Tܕ/ ce/k��4HļsՀv��_�lE�eM�M��u~W,��t/��?���9o0���tf��;g/
�,���g3���:,�
{k�3�3�J��;����(3X'$y+��i"�����$+ܻ'�+���dW�A�M�� p��뿻kY/��g$C����尣�� �<gj���U��4���f�Dr�������� >��������đ������.���u��/4
�eh��/��~~{~H��C�q|�W	ϰ�����!D�,�������s�_�X1����!LZM+�]	`P(2ܟzMV�R)q�ZU+�������ɦc����P��,��L�5�f�m�.&K۱[����;}������׳h��X�)��>E}[f$�"Le��T����ɾaR�zQ�Z�!�8�� ��Ğ��V|5��=9}���ztn�;v=�������B!��zP��v+f��I�$���K���{�fx��yD�>;\�n�!�F��������0��p$�*�CV��bVN�/3~L��r�S��5� Io�e�g�Nꣷ�q`������\��nWj��e������H�m.����=R��k�y"��SE֩YD���anhF�㳄Ԟ~�C�q�0�R���*���w�:�3�NƋ�����*A��
�*sN�\�N�-��^�'��GIK-s�S��~kN�V�R����'&����lF�Xirˉ;�54�٤>�mv</�h�䕠s�����΁K�,�8#���-b�"`3��e����-9�<��[��w^Ç��3��|���Vx��`�+	m���BN��/UGzz���U =����D����J�|���x����m�ݏB��a���/}�)����u�7�j�@}�����hv^?�+�'*��Z�ڊ�m���'-�Z0�r��c׆u�;��,7"a4<e� /M�������g�K��Bi@��[��o�
4��l#�+��%k��Zr>�O�T��"ţ��_5do�q'�6a_�"�+�A��>G�R��5��֋3r��*	�Q���b9|eŖ7{�)��pt���Bi� �>�P0 ��������=�ҡ[�<n1�"D�E2?�񖰦�L�Q���XG����B�1xȕ21���'�c��\���-�?S�x��#j�f����ѿQ�`�]��EC�?��OA+Q�٘���.}�4;�����	�<$|���秃��T]f1�%�ǧ��?�7�`��D�\���	x��ؐ�J�,��}ɷ�u_B�N�@���ϧDG�Q�&�P�L��r���f�6�sɈ�ߢPI���b_oz�"J��5�l&������**t��g��a��M�Z�[B�b󒒜�:���m�0�J�1|c4JZ�j>��Z<oIzA��u��o3O6�q�?�����즭L��L\��ٌk��Ps5��}��ߡ�c�|KN�\¯+w���C�z��B�� z�_���񚀧����%?�g�k̓�>7��S�兏V�56�qS���L۴����K9J�;�:�Z�����++�uZ�Jث Y�Yw��X�L+i@��,񃘟����KO1(s�<[�^�IZ�>V���@S|2���ؿ��{��exY�f~�&eұ0X�����~��j=/ͫ-�����G�'���I6�'vl$	��=�߽Pa�SB��(u�6���䆝Ki)s������u�5R_Nj�'{�E��]�B��!�W��Χ%%l)�x�׳a�f��->�B������ƬKSvV��� e{
�7¼A?lH�KJKb��8䶸����߿�4_4�!˝eNr|�|�3n	G�
��R�AC�@<���㌰�Ȫӊ����Ds���a�Ǣ-={��`����H�^���ͱ���_�V�-�GS��E涼h�ޣI<k,Os0	�4�
�7Խ���<�J"�4���˻z�`cA,<l���f�'�am���ّu���=�rQ��n{��ZI�أ�]"o4�~Nb?+�u�
,Bx�N�0zhd���&�]u��"��el�-�^䯱!4���V2n�K���g�d�t�k���ӿ��P��fJ|��\��U��4~o�����tYń��+d��w�R�D����[�)͡]]�n�Oa�Φ����c�g��Qɀ��'=P}|�'i.�Nˆ���(��@�g~t?���7&��h�j���68.�b�N/ݳ�?�aJ����L�KSqJ�~����\<3�#�\����l ����綘㹃�m����O�R�����5!��gVo �q�O �A��X��F�&��Y~��j�Kf�al�`�Dg�a?�_I �u���$����ƻ[�ձJcH����K^�l����^��Bv�<�f}��n�>->�:������Y���7Z��?_���Z�#��~T�b�P��]�%�����4 (���,�)G��x��<��k μ�ǀ#���)��"�&0+��~9 Hg�9����8���x��2��Q�Z|3�m1z�{�R�ّ`�X1���9o5������ñ���#�<�N^n*�W:�.�����ǵO���^|���'H�E`6Yۂk��g
�~���U|����'" �oOTBC(�S���0�Q.^�8�-gM��"����/���kݮ-�q����s�����^�@�7�l-$�����Z#ՙ����W��g�Wa����Q5�Ԝ8#�+
��GP�yL]h��F>0�(R\v��^�ݷ{�D�Ot�8E�dK
zy�x���go��œ(u��EY${y�\�L|/���u������3c�9<N�x�X��Ӿ����O��d;V��%]_��|�u���D����'�,�޵$���3�5�ė�K6�;VYwc_\��ta�'
0�h����(�S2/���=�}����ѾR��ì��d�/'�ЁQY�1���}��%:�&�qs	r����	4�G'���^��`��RX�԰�ܲ�*�䱃N���W�DYGN��(������@���K���~|����O�iɅ �i��i��i��,��;R���Q"޿�w�#��}���;fޫ&�[��lZ���O�'����e�nA~�v�b��/�8�Ǣ�Ðw�CZ����1t�*S�e�jy�_����b�͒�-��O�rA�'�O��Se_�.1��~c7�R��:�70������G.�����W�~��@(�क़���
蚸I��Hp�ѳV���L���ԙ�����J�x�z!}α��͎�s��Zz�1����]��a�Q�d����������P���#]��N��^����^����I$�N{�[��������b��48��TW�yI������'����-�y-� �d��MG���P���X�Nw�.��w# ��f��Ƿ�{������,|ݦ�=Y����-WD�"RC��h$~ꪙ�����58`+�a,�E����I�i+�E�^<��6�E2�ᒑ����|��O�lz���W����(S8scb�3�'V�ڼ���NjtN��'�4ɪ�ܶu�y�}�e-2� I\T�KT�9&2��8P���T }޽�Eem5�B��AS��F�)!G�e[q�I�T�E�kX����mm~X�뢉Mb=s��=1�I�4g߽bz�����t�����.�f�}�
���X��4g2��;G���N����v�U�k8�u�W�zE���O-O�C4Cqv�C��b�C�'H�D,~�v;��� *Iѳ���q�ؘ'�k���93*�P�b��&��W I���t�nG���6�1�<��0�il���&�G0b|��)�u ��Q����������.�T�E���tD{ݼ�$��"�,���^�68oH�ڢH.G�_CC
��`��+{#9r��eސ或o�F�[.��q��V�JXZud��>q����#{�L�T`Fy��+�^�[0�WRF��;E+a��s@�Yc���@_ҽ�f �>Ћ� ڛ����Ԯz�8D3���:�-��3jmR�L���7�S��?3��ؤw�}��iMI��Ii�zǨo�6��/� �x��<����D�7�k6��@A[mT��̆v�[���sR�V���W�BIE�fR2��K�����>O&�{�u�[:��<�`��ŁA}�����1� gՠ �ջt�����7�K�G��%*�SM�~1��P5���[8�d����n �5q�;@L�L�P\ƩZK �I�i�K�8i�;�Lww�H��:��s�������Z'�w�͞f("w�e ����{ ��ؼ:ۮ��\Lh�����MYn�hx�K�u�W��e�8βϓ9�ځ��?u��o���l�Wǌ��:|)`����Ҵ}�:]�]ܸ*�+T��TV�K��e�C��r5�<-�x����e�P�g�x��w�U�w�[�jk��1�����o�XnÚo	M/��E���%x`T��C�o�=�mQ��ʃg�(��RQ�ׇ���^r��L�gU{
R>m���W1`���š�E�.�1'��#-i��sO��oءD�p���_�*_�!�vm�t��k~�Y������{�x���T:;�c���a����c[w�TM8h��r����yY��x�-���G7��G	��53���?�Me�A�j������H��Z8ۣ M�iC�h�ϏƯ���?铏����zX�Q��\�|��*k���8/SS�`zb?c:�}'t!�(�d����Sؙ:�\Z5�-���ۏ4�"W�����5E2���w˳�o���T�u�NQA�P�m@[��Ī�@�yS���t�7�%<>�F�v����[��KZ�[Su�����d����=Ee"^�l�m���c�3X��z����{�:0���BW. �x��$Z
c�#�c\��Υk����Ѩ/�_~�m����_M�/}�߷#wwٕ����$	��+4��D㧪��#�}d��	?l-$�Ukݛ���T����z,��1�ͫsb��N¼�pBgjsT0���-8�1/�\�xǏ���yF�:}V��yIY��´[}�ofOH%�Z��-_�?k��s���À���@쳐��X���L�i�̞#��;�t�!D��[|]��|�)��/�|��/�#s�ķ(0v��ܼ�I�k� ��s�B��8p���q�J�g�븱�H7yo�{���m�{�N�d�����)w�&�<l����3G��q�K��#]'����/���F�#H�S�	|���y;�ퟶ���|f���*ʆ/U��(��H#��Ȣ5@�����նc�������*������&�y@^���Y#	�8|�uьGan2�}��ԍ�z�a%Ѹ4Z�N٭:е��K�}
t>��ٝ���Ǌ�ё-uK ��MQ��}�㴌�}�����=�Uy������܆�[ڵs��ҷ6�"&n?�����J]{w�;�U�|#�Ϡ�?�$�3��FH�b6E=�Z��y���*��5Y`�fD[�CNS5�!�	�ʴ����j�M� �*��$����k��d��� C"�B7wT�6�}=����G�&ո���T���ei� �߻. ����y6�������^E�\��g������]��-��h,�d!	��;�[a���P��ӠV=	2@9�e:(��֞�ԥ���F<lG��<hK�&���tϛ����W]��G$��J���a��z��ETF�|����ҳW�D���r���~���nL�v���r� ���ڣ�<���2�k�m}�Ik�`������z�}/ _��}�5���7�%o���d]�i���E8�&\�d?F�����}0QR������������hXF�1)3��=mo�G{�����}��-,i0���)�P��A��v����}y(Y�
S"���o4d��>���	��T.kpa臢-�
��h���z��i�-��7��ڗ"���|K�7!�ӳ���a�ΧP�j�{�D��7�a	��C�c�bB0DC�������5���Xl=��������p�����n^��>�]�(�U`��l����,X3�����1HM�O��#($>�����$�l�d'��d���^�/��R׬�oGsm`5 k����wmԻ������ϟ_�Ar� _�6-��ύ���&���{����?����>鑏UqJ˒rϽ㒩���nΏ�Go��yv�-��
��|MOϴڔ�N��X�����/l�	}g~s�pe�������- ��K�B��/���Yx�=�Ƃ��z6�ȹD��С�;ۛ9=O��"�+k�c�PSn7-j]陸�S�����(����և��Ҟ�^����w�����tǀ����m��S?w���o�,�^��/���鄲K�m�� )4��1�PQ����EJ�T$%�E%�:����cH	E�N��nZJ@Z@bH�a I���_�����Z,�;�8g�}���2�Bû�b������3+�@v�:J2�Ƭ�0��V A��O�/NXch�N�˻�����m��؛�{<��P)���������
W��O�4Rz'�����Ĳ�*|?aEN,Y�c�r\j=���a#�6���mH�1\��~|&���|�|�LUi�e��PZ�&;�/�~�'#�+2C�}��J%��k�JSA��'[kU����E˥O=�K~�H��nn�ں�7�*3�{k��N�b�[T;�F|&d�ǹJ��_7���ȏ({�X��"X���e�>��m�K�U�J�o��F� [���Q���,�Q��g����s~W�!���>�E.,����S�L$�C� �N�VuQ��6�E���$��W���.J�9���:��	%���N�A�|ؑ�*�٬t~�[�u y�Z�����1�I���Ҕ��')�gy���}CTc����t�	;ѷ�@2:b��er["�2fF}d�8O�
D�	*0艿�s�lR�������&�*�͓ͱ'�*��W(�} �.<�^T[#��1�+�ĩk��)�K#����3l��m��-���]*I�rk��wՍ|>5��5��[����xaTNsu4[r�{~���u��NQ��91�%���Ν̷sm��?N
AI0:aږhV	g-��R�,��G�Z��:�I�D��s�s]����g��O�|Ƴe�9P��(.̥ɽy۠��.I���j,2%��5�;qxLs���*�Fk�rZ���3�2�%t3�h���^��	�֜�D��Y6|�������+�I�|֘v֠��2���^����Zʟ,Q����!�GN
9T��ms�fZ�Zw�=�1��e�YZ%�4M}7jH��~.ϲjL��"D\�Ӑ��ᷚ�b�+��	,اDÄq �idR�޽�rW-d�3�v�������WKSJr,B�d"�??*� ��w��2D�	����bjo��zCY��]��$�C�˓�����OQB-��>;eP�<��%>���]��-#���#��=Z׬F��Ȝ�s�3�3
zS�|A����&� �ٛŅP)���48(	`�cqM���wI�	�1�K��4_�ǜu�m��������v�P��Ѽ��g�n0&�f/������'�1�=7�����̈́�+3�4��	�i%�@y�6����]ňy�m��5�Pj�v�gy�
5�7r����V�G�O����\�쓝m�8����a��nac8\�	��AEw^��'�P9����A4��(�Z.L�T�/�[H�ɖ]Fڲ�D��~�a�����ߦ���!�3���d�`6"�4�X�����j�N��A���9<rr�B�N�Vb��Id!�c9�\<����B�N4P�� �:����w�!�A��U03�G��4
�(&��!�0�9 ����˼�cI&�)pU��\�喾�"ԋ��Ù��������/��X#���O��\������ϲ4wl[t�����Z�8�:����򊍝��d��jźl[�{a:o�Yɓ����/T���[�ᒭ���PV�~WZ�5{:g�핒V<�l��y؎���q��$Yx91��#�����봡36��q�z��a)��P�b��qP7E�O�1��|���ڸ���"�M��zr�J��O0��UV�&	گ����AO���)ٮI:��g9�?��qX;2�| w^oTE���6u�M�\P�f�FjO���N�&^��M|٨ �gs�0��î@�	_���g�^�ݮ�b]��6߷�����̻��Vp\GȘ�Ud������������$�j*A����mϗq\�m:rb��@7���.�ԟ��y��܆�1��Óղ�Z�L�z2�2i#����p��M���J�Y �.�`�OQ�.YjR;�xч�bL���M3ʡ"�n~B�2��R��)��V(�9�:p\m�A�8Ig��l��Đo~��f���T��j^�����*߂��Jl��٪w|×~�r=^4���1��Jj�\%�*`�/Iq�@��o�J������X���>�ri=��Di2���Lݹ�O;8J2��a7��̌鎽F��}�Z�ן����z�����˪��6��!yQW�ѡ^��ά�nK���2�$c�����M5D����7I}��lm��ق4���$s*0L(��z�>�j�C�����uגH�`�#KWZ�R��ړ��,�,f���_�͑�r����wv�a����$Hmuw2���A&O`�gcf}!��AÔ���T��~�X��Z& ��qn^�x����Rk�&\5Ae����!r�`⺂?�i�7��P�$���橲��µ�y�0Ws.N����/̷�O�h���8�%>�o��ç��)dq:K�&|ឺ�n7�ioI���o�E���8�?�P|\~���77|���isvP���Td��l�6<���jX�\!�S�+"�U@pJC��Ug��[�ٓ����۩h�zVY,�Sd&$e�e~��_?N��ۤ����V�g�W���d�>�(8���8��ˤ	�3�N4d&*��p �N��w/��0��[��$�, �k>Zb)��;-oN׎p:��ZvNP�"RwV+����8��q�0Ԛk�K��j�뻣�Q?���e�I�=��oө��0�\$M,�<C��Cp3d�?��t�"�8�a�O����%{��G
�M�[�Q��l����iمX�Y����^VLI)���n��a��x�IL�,�	���km>��>�o]�m�����֞���;����SX$���#�6Ȁ��^���Y�&9G��e%%u����;?	�wmdH<��V�Ot4j�b�
��K�b8I�J0��l��@D�w;�8��ET[�/R"��r�9sr�.�+�7C�uO�FŤ$�6�r+W���M,1��'1�®�UT����#/��/4]���'[��f|������ĜJ5�;�y�W�ae�; p������t{{i��B:��l֖W���*+�#�;��O(:xy�.�W ��2��u����g<��և�f.�6J�-���&����zT���"���ʬ�4�-y�؝U��(x)ى�%����o�=ϟ�.��n�(	�MQ꺶��hTܞj��_��b)�z�|"�ɲ�Ѡl�t�v��|ͧ>ؖ��xp����wLJD۔S`��M��Pf2jTy�>ZI5�5��d<[H�w��3�q�͏P$�Rqm?ܮ"��;�}0���> ���h��z�Bb���/.�����|�3O�3��1�k%H�f�n4��}���I3,v��D�!����DcRև���EI����<U����cˠ	}����QbQ�裍�$4(��8@�>ӣQ�fM�.�#`����a��w-pJ��k�c��A����"]Z_��#Ϫ_��d^[��q�!��r��RyA5�̬�����.!`f�tW����n�Z�� ��݁�N�������?�ղ�,u�MKʼR�m�hQ�՞g����@�����l����͟vs���j�v��_*����v�j��\��f���Z}�a�p�n�S�������x/�l310U������9�J0o�i�[�����c���^.���{��N9���>/rx#�VKP�;A(��u�g������7�P�d�O ���+�`��4��2�� xv��-�؞�Ư�i�x;��m���{ŠYUvi�>�=x�2.g��6�n�n�����6",T���a�����(:�F�q�I:�)ie�d'�����6'��.��u,f�~�<������.�v�������оq��}��Ӫ��0���~S$p�C˥˓܆ER<Zm��2�3�� 'V��W� _��1����f���k,Fv3�o�������a�/j�>���Mx����=�x���HҔK<�p��ݰ����~�����*[�v��|?>��[��U���#w�[p%IBvߕ�t󼺮5=�a�9w�o�L�[ވ�i�\�V]�9��*?7�#���8[�z��7`p�m�x�r �s|[��؇�E�i�D˷2�D@k	l$>����EY�SQ�����)��|I y���f��|�>`,��|wW�0U��׈� $[ˣI����wH֩�vw՞��3�E���^��B���#�;-n'_�Z�KD$�����{����u�u1���r�Yp$)B��˼"D�W�t
+�j�$��'�a�����`����s�$�0��!�P`w�YF�,`��9���U�?��M�p����zT"H\��g���f���\��O���N�2����T6Ӡ�g>���(�G�$|)&$���]��:��8/p���%�W^��b����菟bCwd��L~b�p�q��?e��T�C�e����_x&�"j3q��._��x@��:��)\���f�+��#�BZ�F�g�� ݏ�?�c��44�ug�aNL��=Ӌ�}��r����/h�T�VWV���t�V8�A�n ���X8���k�$�&O�<s1������w�v��F���7�A>��6�]�d��$���)JϬ&���雾��#��jJ�ȑ����� J�w1(� Ȃҹ�r��[JtJ*�ޓ�c��Tа`H���zr�bG������[f��c:�U����%�����4��S�nՌ>�X���y\=��$����Fz+��oo1Mr���0=W�m��)��x�k�&�����H�*�GL(!��EI������6ma�ک|�y�}��,�I��mZ	�Q�,�x�5��e�l�~���0�4c�K}�RB�_Zm}��}�`O�y�rK���%�b�\F=o�L�Z�F��qaޢA���B��()�TƌZٱi2M2qj,��F�
��'f�'����eƼ�S*������� �On/m�w����X��
�*����o�oLj��?��r�H �<�ƒ��>v��,��:h�)M��D��KCb�vM��o+�,I�����D�o%�<�D)�l��2���z�œ��w�I2��ZO��&���l�U��#m��_�H��"){���?�[9L�<��㻎��_����Wz��[�%"߷2 �;���Q�un�$��~�-��Y"�=�� ��r����~}�"�q���V��|��.���>'���ͽ� ����ڛ1��y�#:Cߋ-7YqW�艁M:!w�#�I:�O�Q��s�tޅ�*��Ґ5_�ww�0�D�.rԓb�{�����!s�
ǧ�'m
iz�;`u�)=l��񧶧,�/���UOѼ
�a~����a��1������Y�����C3�(E�Wƙ�r�T����N�˜I��ҟ�H�`ULj���D������GM�z���El�a��F2��Q��6��|��e�Z��N̹0�{f����f�w�O� ��M��s`�<���>�~ Lר�X������w������r�<�Pe�3l7�Ӻ������F��̗�J�r��v�K�[_���m3EZt�%�6Ƹ�Ckw�&�k�����nWL��:.(����,�[�|��lVakQ�]`����`�
O���H	nt��X�C�b15QFȠ$4�p��iK�CJ����Ȓ�������Q�F���W;�*S�Z\�hs��T���LYo��lּ�t��Q�𖍂4Ý���ґͧ��S���r���7V1)R�����{O�8nثv��D�n`�_�)ܳ׃`�l=4.�#Z*�3����s����0F��ܓ=�0�؝����/�v&�}�K)3;�Bq��Ӡ<�+ ��h����;J��$b���˓���[M�N�xtg&s<����j���H�����P��E�ͷW[(	';Y09hcj����@�IP�l�&�g���o�5T�#~�a��崙2o��T���3�޳?�����9A���Y����+f�z�W�5��Rn^?5�ᥚ։��_4��Fj��N�Vڋ{u�����R�H2��n�O\��6EF� ��Tiz>w����11����S��eM˓�-��6��x��ּ�fan��ǀn���#���11�Fa�b�4�����"<\=z'��&�~����a��/,`�>�A�)7L�ڇ�6���b����ɏC�J�͆��4��*u�bӋ�����wQj�GYwa�	$?V�a T1���Y :�r�U�O�0UZ�62 �S3�(���JV��!�d� L@y=���` �%��Ȧ�^e�oL5���UK%b�6Yq�q��\K��֭L{�ԍ�Ls�R�)��W�T��}��˕
�jl�h�m�������ݵ����f�d&� v9���WS�	��|������*��@��?n�{�*���T�Sk�W����4�isT��h�+�0�l���2.`l��H�t��z�5�|�|LBg.�lMs���V�\�j�	���%>c`�
f"/��9W���p�g�� �A�6<���aD̦P�A��u�_�&3�A
�$�F?|�H�NnGn�6�� �7���<�6��:5༠0>��_	�����'�B��C%� hB��5~�r�؛����%�!��eW�_�� b}}cסuFyr�c��,�*]F��m�La��x�����:�;��!�ڗ���p$.�zI�^��a�L̤>KM��������6#�U�K�V����[o��T��rU�EXE�ߑ�Ag=U��<'��z��]�Zm�]�H�>�IN:����t��%�� �p�<4��;Tu9��1�`TzmJ���6��i`��������7���I���;ꉏ���Y/uDCa5F�<�UK�G%��� MZm|�����q�w��ٴ˸�����n��$��3�'' С���!���+��U��<r�T���x��js���j0��<	��0�0�k"�� c�F}�vǉ�倌���-2�����~��w�S���f�Ϋ/�]�������4�\��ff����U+lGc�*�?a�i�k&q���s�9)����4���M�Ta�0� �f�2��B�[��o=1d���jR5dlj���\9���)l@��Ҩ�6$���Z�v�\��v�̀"����Īt�NB�͒�,�vz�>�LоEf��{h�!�&\r��4�|��a�@�� W��BWM�e���e�'�ڄ����c���ϧ����W�١�z]�@/�H��>���ݔ�e��#Ű
,�"�<������w�I�(@<i�#�횐��R�k�m4^�~˫a���w��c�׽s���p����B��e��%�t֟2\�a1y���T��ݩ�ds�M5x��*��G�=��OW���~�HO�S�~���p�z�\��a�Y�����G�Mߠ�0�07��p��E?b���¥9y)�?�E�HɅ�ȁ�����]p�/�o���s��^��c���y%ܲ�r�3�fAQ�|��?Z��R�9��A&�ˮ�i��xn.X��幢Y��A	x��;8V�#��l�3�z �i�&�e�Xr��_y~ф���U"5t����4S��=C��/2:�l�{d:���؞�?4�?ϯ�ez��Q����bcZ�<���T��pS	�hll!�WAr&�c�	��;�_���1�i6S��J{��w|}`��oqD
R�Y�Eq��(e��TR��d_��X憗���#�����6�|^��O���ڞ��		1���������=�����SI<������x!���%e��Oa崯��_1��"�`����zv2�����?����	�zJD>.��2ZM�O��vRHCƽ���"�I�c����\s������
�[�_�ҩ2�t󁍞njg�(�܏O�a��EF��O�MxP��z�}�7�q�����5?�-�R���k����o�)\�V���ly��=~�P�aQ�c���&�<uU�U��f+��l��n��v�9�`!�E�q�Ⱥ�:�8+nBN+3?b'�¿�՗]L:�=��}2��F�|,�rE�ʰ���1�e���i��L,K�<���w�FV������|R���"������/�W�L��LY�K�&�G��,H.��q� |]h�ev�,���2Tȑ�T���C��$��z��H9��Lf�[�!���<�����H͵�l���������:�����ƫ�I�K_��<G2Dr𑋛ȅ]��w�.��/�k���b��иͼ����O�d�Nry���OsT�`��A;Li�U$
�6���o�5��v �8wm�"���q�m�z�M���L��~�o��w#~����>�]�P�ć_˼�M_c=�!\����Z�#=ܞ��h��3�<�ě����f=��b�v�������^����5k��2���0�����ï�$`�� F�3�+N����.pP�E_�Fے����m��\��ao�nN����$u�?_{h���v����+U�(:��C<���E��t�3��`������K<�X|-y:N�j�-G��ɽR�DL:GLv��`�����ΰ��$\Ea�s�p���5z�N�g�������
I)w�oEgJ�"M����k�Xߍz�{)��@ĺ�y�%!��l����i1;�������kB�,j�?k.%��\F7Ń�=�g�PT\�E4��i5q�����{A"�nz �-1EO7.1Et��'L��FP.�"j���[�@^I��S�GsMr�j
;������L��n̳�����ޜ�2s�ޥ�	���a�	�gV����tե���^k�=ޜ�*Ϣ���ld�_zp�b��='*͜F���B!|�i�F���1i�m���1�k�n�c��җa5�o���LI�	�=6^����V;��o]�ٍi"��kӰF��)��Bs8�C�]u�L��9�K���)�yw-�!s`#D����rw������2L�Y����\u �=C�T��ȅΥ�K���2�?iƭ1�H�v2Nr 6���Q��?% P3U��v�+6�dF?`���&��{�ãH���u�8��A(L� �ܚGv��Z����H���?YA̧I�e5%4��s�}��,]���	΍ڈ�w2ة�ša|g#�+5��&�������LJg��8:���n���/�"1�n��*�Ŋa0�lww;��=֤�i?k�a��UK���B�FZnyŎE����E�L��Lӧ���^2E�:�H��R����t��L���"�v�EË���:(��of�YЌ�,�e.:)"��(��n�&�N����t7������n�ǖ�	=G�T1�*pʕ�]�s�jn��@��]���jG�iyu;�gq ��e����n ��T��r�C[�8�؇lb�f�6�tB��j5noY�3�+8���xcuʹ���#^����pn4��M
{w��E_8�4�? ��@ƽ�'��=��d���_����P˕���K��q�&?x�:�I�=��5k[����!�@{�إJ�S�JF��I,�����A�%�o���D����t���P����j`Q�M�Ƹ_��
� #�-@m.a�ED�{U?��Q��m��JB�L=�d9�Z(���
�+:�3e�����Y�M|�W�ޮk�*P�U;����N�Z�׶Eы ���o�HM��ͷ����Ƒ:Ԁ�\7�:=8_�̈́���	�� X�^��Q���_�m�+~��-:���is#)M������0:�J�����T�� ��mSk R�A�/�\�_8g�v=y&��RR��5կ���D��/3'0�/�]Ӷ@���&�`$%O
��ϳ�o�f�
���[R�	��h@B�wɃ{�,�������oH�?�*:T��y9d��糇/�?<7����>�^؉���ZfGg_�t�W����_��!�����Wr'���l�������y�	����!1��:��,e�ю�~w3EHw2�p�ձk�m����'_"�]�� Q�� a&�(@S!���url�Mn�:҆��o�|�X"��u�=g�������u��y�U��>MC���Pq�'�s��	�\���>�ք�:`��ӎ:-i���Ma��z�)���j��>%BA��F�+-��r��4M�=B:�:;ܾNfQ(���BO����DWa��%�	��7: #�8���6;h��!�����;�zF&�ϯ��ܛc8�ѼOp�Z?mh�_���l�J�CE!rU�@�Oc(���Ƕۯb�ޅ9}�뛲R�#Et�>u�&vт��=9�|�Q+��n���-�[\�����E_�Ŕ�g��Wi�d��EV���k�A2��)��L2���#;>��1v��LR��!��N;����<�WW�оi�A��{g4ל���}��K�G�J�T�j."��Cĭ0��L�~�+�E};�Q$چ�nڳۼ� �~�S��sWԛ�v~.�_�L�]}��s���fa�0ػ�U|�
���)�^�A��ea�y��E�6��|�@r�ޘ.��>��fbj}�I�{_��H�>zz�,u?,W^ڇ8���<�;d�gƅ4�6Z[�#�z�V)����]�r�R��5~�le�T�٪A�0W���Y�L��T\D�=;��gyW�̍ޮ�7��2��u�PEI��}=�)�)�`d2�dO��d�j��V��U�����OZƩmȰ��QW?���Ih�ݲ������?��x�*�Oh�,��JEӉEe�����ĕ�&�L����l7�B�|��E��Z8�1��L=�JY�e��cܭ
.a�1.�}D���h��<L�W���ə�@W�U��uyA���i�5T�aN�˃�&�����VG����*w�2b̒��we�-�GÇv�zn�j2�=/�{zWx���5��N�IB�oOf�w�٨�J��	�U���q�Hb�ԃ�!�j�o�.��V����qFv_6"
��?>b���g3~8f u�#F����g��/�=׏=�w# ���i��i��d�l��As������C?��U�:�����~����F�	]��_�\F��y&�Kx2�����3Śi��py-ə��7��Y>�y�1^	yAm��ƹy��EG���Y��Q�/By7b���Zt5��%-��Ӵ��J���[)����y�����������4�M��eJ-耫F6?z������^�v���^�{�L��vm��M���3�ӧG���ʇ��Ȥ�w9$#�*z=�̍���L���o��Fy8��s_V�V6�%��@�=l� �,a���24���������\g6D���y�������ڗ6E�h,�Ψ��&1�}7b.�iOGj��,��PZu;}*����{�<0��=x����!��7��~���Æ�5{n���o��$��ظ��d�vV;�i�M�����hx�n.�i�����5E!zt���D��� �(����"/�n������SNk���ϚvU�bԝ�v>��)B~HC�E�"}%0pYj���Q���a���^}�ٸ����}�|9^��J��׉0��>���;�������Q�n�tCbz�:�[���Wڵ6��,�g�1������i���ʸ��$���n�&�`��:<�^�[�L<O�SY��T��pp>��_�E?l<�����l�?� d�6�.!񓥀�����>H	�������j�7����ǒK�1٪�B?��*�V;}؀]`�|)<�;��3������>~/v�2�+�n�o<c��	p��QVW@��\!aa*�L~#T��4t'¹� ��u�ћnm�yol{��)�#t �dں�F��������7�����r.޷�8���E}�+r+�p���aސ���d
�o%V�[�+s�$�M��#��4��D��������M&�Ha�S`cS�>�_ 
�IK���N���>�$��}�mwQ{��u^��	<��Z��&<�os*74zq�N=��pՠo������9��7����5ɖ���ڳapحH.��|���?=�����v9J ��U�{cV�\�^�4�cC�����ݪ�}+�/���1��I���m����@���Ta�(�`6xb�q� ��)����̄z�/���=	��G��j�`³."��&~����"���J7��߀5Y����8���Xy�A˱��A����N\
xӝDn�dbXT��m�V:3Us�7$�TQ5B��x��<�o�Tb���G��a[�n`�|-����|����V��r���Yu��|�9���w�&e�g�[�0p��9�|�s��_Q4�0�T�О`�WU ��P~�&�~#�bcbm,�A���}����ٓf�a��?փ�Ε4Qp�(�Ь㇊���R�ذ�7���c�r��R�d|a+,�iÚ�����h�l#�¥@��|�@lm��\��Ll'��?"ur�;��E
'��x��X��C�鿡[��ו�ƾ
�a6���z�� Bł[[cb�h0�;�+8�<4�_���1[V#�HW�����\�awf�o;��re[����/�J�lՋB��ҵ\	w{5��E���f��4M�X�c�o�\��'iH'M��p1����@��W(Ŭ.�V�b���Q`([��/�jx�y�嗹�SC���b�=K8���f�ьN��R4
�`���U��NBρv�P�m�z;zUȶ����숏�z>T�=9���8�¼T�2���?��n�'L����Cu��<j����R�l�c����F: 0Ա�F��̍�l M�S��L�7R�Շ1S_��ex��<a����A���GBV�{�����<��ĕ6B�K��-��R��3)�ŷ�۟��,Ƀ�J`.��\#�kz��j���eN|��
έ	yS>�����Κ-�3���gh5��)�9qʛ���������ˑ'`�X�����&MbeMZ�z ���\����lh{�s��MF�*+G7�7������D@���2�g20w�Xod��)�h��b~�Ø�B�Y*�-��2Iڡu��;���Vt���Y�(��@�L�f�����ZpNr��Ç���V�Ig]�jV,��c��~��ޟH=��������U�^4PD�&��d�s�e�o/��3hX����%�ދ}x �bht7J�F��*oɅ��T?���G�K�"ҋb,�R�$j�E����Л�!��Ոi�=�M���YV�ڋ��>�s�W����h�悄��E+6xQ!��}��L�����E�kg�r�;��kE -� W�Dw=a��N��Q��c�!V���Ӓ2�|�la%MF14�0lz�Ј�6�YG���'�H����l�0XHr�m�S�Mj�!��^~��MFf�39���ظ<����g��I�("�A���s�&x�D~t�&	�O IE�������R��b|6J}��Z�V�f�۽Ql܅���/�C�m'�FP��e:et,����V�a\�-
H�rp�A`Q�m�d����(��XD�o$Od5O0U�,���k}Ƀs���sko��99���� ���y�Ǘy���[�ϭ_�zӘ�FC|���c���r��gMl�N�]Pq�RF4��o/�꙱�:
���(pg'�2�BH��x�Ɠ�4���V�n���9h�T4ʉ��w���׎k��!t/�S8�M#����}qAseR�=]�7Ɩ��H#hJ}�i�#;Rk�h�7WB���`Pu�G�J�E|[&���v���ڼ���뫑CIc2�[ZZ������%�����-�r#]�!/���X��j��,Gy��� ���+���	�o`AK|^'�:���g�ﻎՄ��J .v �\��s{�_�����6<#B��8���_�̶jt��E��].�z�Gb��s��凴T!���)�B?�n��H~ֽ�� =�p�B�b�BK��\��%�;��֯ ���Ϧ�B_����_E@mcyJ�fj?"�F1��A�A4��V-�X)�w2���Z]��J&���8�B��X&��z���4H��Sb�&>W'9��+��b
�Y/1��nzsv��ȿ)/�f��Ü��ߥ�ʛ� b	A$�RN�����ۏ��9+5��ԁzj�P��8�Y�LJǠ�)��<�J~<lK�Q6@q	]ua��v�u
����z���>oO��]�?wg����
B�I���b�©1�7�b���f~&O.}��*c(�$ާ!ĩ8i "m7T��K� ��q���Bct��R���D����dJ�p>������;���R�̕_b΅A����y?P,*�O��+��^cË�i(%�m��i�v��H]�Ѵ�"H_7��$Jй;���X�|�Q(������@��Cnk�j�s��L�9O�����3�SG�h�VV�q�E~���T�D��$�B�'��[ �T��G�GWIx�T[$Ƃ��wK�R)~����=~B�A�
��ۨ�����]MS�m̱J��[�ß������s�}aX�vt��F��>�	QS���,���u��g��[�ߝ&od���f��~�W$�L=b(6;
�R�hfQ��ג�b��VvŔ��r��
���Y+�|m��=l�B����e��w��cğ���ɨ��|��Z'�����+���P���Qj jb���+��@�Gu%���7����?�x���l�#���xzC�𣍕W�/G� �;rd8pn����c�����䋩�j�Uy��K&v��������o{�:�{�<�hq���Q,�;��\A����X۟��_M�,�J�����?sVTN��Qd��\���#�%,����db0�T̟>Z�JlH֕�X�&�Ҡ�BE�%��?��	��f��>@-�N�I
��[IFlp���kh�X�f����ۆA�����#d����8���H�T���gEy����c-D�����	w�T�"�agc�`�<�0��j��h�5���<��ˏϜ�kF�ۡe���p,�e�G����I+�yl�k�柑 �����g�����/�s�}��T#��.��GE�O��`��į��e�F��1�֌p"��Nl���7��Dx�w�j+��`��Q覐�l�X]�'�Go(�+o�<����%x�h?���<�YՠMZN�9Š�9�;ܷ8�)�WE�9\��pAu�P|�l���?z�yu��FP���n��ׁ��;XK��OZ��ip�����s��f0��:a����$���{(G��}�u|$�˿҃����{������#h�6֛`-��u�N>~�[Tv���A�t�l%�������E٨rB��ZS�������g�1p��Σ��T����訤�9A�G�N��ȎQ� �#�� �<$��}	ƴ�i�پ۽�3M+�w�"�x���l����|~~��e�:J{sG��4R�du�Հ�~��";����)e�2��Q��@�r}�>uǐ����1w����G=�u���&�<gg2W2��q{[�ß���¹���#�mV�?2��c=�3ɽ��O�
�q����b�6\���]{y�124A%8r	��**���t�S����۾���jTmnm���9}���Ӥ�Ҁ�S���T�K�!}�|[w�t 	�BL�����44��S�Ό<p|�~�
��7�ȟ�����r��HO�E��y7oq�ȳ�N��%�[4*�`ᣳ�he���Akߥg�����`�H^~���<�ʳ�/�f
h����d9����\�3AA ��ڔ P�x`p	��7�9[KNy1厓�<zsp��la��'M�od�>PQE��p��Go/}3Zug��<LOP��zBˣ.�����t؟4k��_�l�4�5
�j�fo�l�
��X�A+b����g_욺�|��ۓҨ�������!�8x�3C+���]�ჽ��U�'L���!���v�ѥL#�_hn �-����xk	.���ʒ�ң�?�w�]^�j�k��.��8����n���i\�_U�P/s��GQN�d@��A�ord��bx ���7a�����+�k�{$��V������K��?�*��2��`W�w*�F�'��Ծ��Y�ϰ,�A}��Y�*���ᾭ��`#��2��eT4s?��(�)K�&#�ͯoo�-5R{m�髥�8���7�8n�F�$�Z�ܪ�T��K	mu�T����]���mk�#��\[6��?#$�ّ���JTm�#�ԄQ�����R�P�:fhG��wR+�|E��a��.�;�:�>�\�����X{	`��b���y��-��d"\H��O0�M@E����!^��z�{s�4�)���ֈ���SNX�u����,:��5�-�� �r���)��6�������J_�1P�}��4�*�zb�@��y>�@1g0^�͛��xh`F\��#���Ja��U�����,Ln�eaiкO���x#qA���ٿP�Ck�8<��5�3��|���j������C���Qn�5��K��u�W���z��~$��fT�.x4~�ߘIF
#� �:�GexF����T�����:_�=�,z�"!oA��U��#�i+?H��X�B���������UA��1	zR�!���.����z�o�z��K]]�bB6�#4o��w��B�W�<���x�'E4Ъ4��y|�1�y�����k����1�b����t���L��)jN��s�|`�}%`�������/�u��X�2��P��TBe�JM�L��'��}�x��TRK��%GY�[�ě�o�09}6c��u�NשG�X̻3�Ul��eV���T���!�����\>�c��d�hZc�6��O���CZF`9T,ɉ>p�S��7G�J�}����R.�j�Y�$��糰U�ކ����L�XY.��0�� Ы�l4����������|G�'���5��ۗ}e��c� 
��;�m�d�n-��` �mK���p?�:����nj�d��5<́��yOv���������-�jn�� �*������;����/WQ��RU��ޫ��H�A�Nh�G�T zE�4i��"B@z/	E��w���~���y2�̞��^{�I(��O=���yixУvk���QXP�ԸWf�?}Lz�b�s�ս�㞾��ob& `�_<��B�j<x���	"{�9�ny�à�s�~JrjM�Ζ���V���+7���\&�/q���D9������mؘ]%$��r~#T?tM@������jN;π��׾��{.?�P�(��դ�#��[W��gd1����㒼0���	���)��T<}_4#���!WB��X��LC�&����O��N*tCh�n7Z:[]\#�y�O��p}�����Re85N�B��ܗ͵�e�,��6�4�I�;���?��.VKq�ݻ��$T,gdD5b�od#?�r��w���V}o�A�Kg%�6����n��O;��3��L���G�H}��~�4�����̉����`o���&h�+"lw<W�߬T�U�#�$���t�� �m5��n�&��rLk(_'�n��{�#>B�'��~CM�����t�5�gX4�OuUҋ�<��y�ڱ:8z�ߜ�4��j�Է�w2[JR����D����<��
���c`�Ľ��ϣ���t�|��	��5�4���BP��w4���{v�'9����s����5Y,��Ui�H��(���v4��p��FC�Ê<����ľ����ܦ����'*�]8?�sEf�x	�_Qmm�Ѕ)�x�f�)H�oz	���9Y�(*�R&* &_����c-�]}��L�x=�|s�x�%͒�I�eIK�=bP�����o�kz���kDWsZY�����"Z�p|׃)�^`�*�a��x�!P0z�n�;�����te�ZW9	����Ҹ)��!���(���ë���u	"�<�Gv�+��si�-�V7���t����cE�w�I�@^c�!�D���Yrb��zkZ��o�W/d�}��k=%��U��dpV��T�M�L��(��pd
���:�� �$��� �b�@'u��__/�L[���� ��D��2���`�����?���)��~0rm��P8d�)h^�Ͷ$�ڎ�o���&2�ٵ<2N�i���,���AF+G�a��gU����S�-m���x���2|\�j;�y�G~a�r�,�G��$<c_���cCC�*���	F��,����e����(;|f������z�h[03��K����k����Fo��L4��2�Wv�Z�����6?�/벷�AE��u���RA�o(m��S��\�%{sT�p%�mH�$����{��X^:[�(r4r�������7S(=�$G�@����������ƥM,�<rbxIG~rv�#=k��+�"���D|2y��X��t��%��4�,b�csEFs���jC������3Q`���Y�Ӊ��3�	������hl$���I��\�PVШ���!�/W��`���O���ݣ����O�7v�t:���D\�dq���t�$�~F����vF�9�c�~��?��l�h�Ŝ�O�t�sR��>�9��as�5,���%zbP|�i���Y1���]�viL��zmV��\�Έ����]ۺ^�Y�@u�lv�q?*8!u��s>�9X	�^+<X(y��I���<0Wr�Q(��Ö�mV�����M,b��c��(�}����ũ�%�k�lv���%!�D?U�4΅Y���r�����5�$������7���U�?g�X�df����;�m;�|}�dz.JA/����B ���9�f��M�O\FJ�w]��L{~+��U�[�
8��h��
c3���\�ޕٱt,T�f��Q{�+�_��DMρ�%����ܬ�x3�]��?�=pV]XX�zT���TF]��$Rj�G���1��[�ͤ)��`�{s�c��_��3�k�����RX����w���]��[`����h"H`�+�����V�u'��բ���A{C���P�!%��9o{Ô�f���>~�5�}"x%�����*�����6s��|�>���^ۤ`!^{e��q����X�������w���F
��]��=���s ǜgD�]p�\�{JfN�`�ڣ�v�B��SVȈ�5��{�{'n{�7e�0^a������ �9>���AG�8�������Щ��:��F�Zp�j��Z�ǵƒ��K�g8��U�Eڰ��P�Z��KF^y�|�w璜�v��nE����))0��L*F)f�
\D���ϭ7ז�������?]Y�jG��]OuY}LL軣7�Q���qM[��|�*���1#y�s�l��of�������/��xs��t�6�}?�4@��]��tDsA�Z����e��I��`W�e${�n׬��pG��5�шKz�?}W�]��9�~u 
}���,:�X&g�JhD�����j�iQT�u������4���V�&e�פ�<�|��=��xV���x��n{��k�z�<:Y
��>��vq"����ߊn9��=�x�xg,�bʍ�ԾKs��@	+�Eb!Z�H �|�� �Sa&j�.�)6��k����s�v�QF�I����c[2Qm���%���.�x���L�Z�������`�Wy�N_sY���K>:�;����;{8o�c�gB�V�`���Mn�/��>�.d����	��i�춇w��0I�(�8�'zi�(LDS�\�t���n��
q�L�x�f[V�r oMoD-f���$�N��wCE��_�=���c���גA��~��"C{�ֶ��x��n�;
�8ݖ�e��е��X��i��P䝋`�gqz�ۗ@ܱy3���+����b���G\	E?j3M��/��ؒ�X�N���M��$H&sj�)��CI������:��J�E�U;KW?}��"N�K<��#DM�9t\�Q6k���yEy�Pѕ����?r�M��t��Di
v\��ʘ:R<vM�Ρ������>>u7����o�%������
3L��������~�����1��m&13��w�s��mI!I�nMD9�a�q'q���Ω�ß�fឤ�p���u�'lTJ�ns� ��/w�9��*�%;��G�NUR��J僎���\�86���jSK�N"�S����Sow��N��2'<����mL g�z����`9�R�]6�w_���������uFF��8�M����������bɴ��i'C����D�ݺ�T��؃oa:��oVE�|
�jiy�����Xj���]� L�6n�&e��5��?J���W��2�\Jn��	�3@c�6M��X<�hz������T�;�R����Y�P�G��j��z^T�⃟�+Wr=������P���Fr�Ȧ�� �
n�st�<?�?v��"��p���R�F��#eV��	mDW�˳Fl5&�
�t��wY����63Ұ�4l�{Q���:,����,�ꘈ[h��O`9p^i���詷�w�Q���;/kW9����?�o��o�-?���Z��YK9
���w�4�%k���ޅ�b쏵-����8�T�}���ؠs*Ǟ��pk`�`c�Bi�Z�(�Q�M�k��|��ڽ�!�ֽhU�� ��G���e�u��F[��sO�����)�O(a?5��"ʑ3,��J�+�����Y�(݉�e��q���3�y����3�Md�	+6��������$`ˋ�����
��_��X�>�T�,�/3��+0���/ �5j�QKK��77 ^�ċ!����d�ib��������>\U�U����z��~~L�q!�$���bX����ȫb|�W.Y��K��l�V�F� � ,��U#h�iN�+�b�I~�8LւX�=��s1�c�Ε�x3P�8��.�����p�ی������ �5�;M��
�*2��LWW��d�9?Ǯ���>hY��2�E�N�H�q~d����y�y�k�K�gE����#b� M��6Y�	��HhsXJ^bwI-*�y�T����G79�� �{� 5y�в�#�-�d�0��c��ݳq��5Z���>I��E�I��Rp1�d�k��?�[�]D9'��$��=P4�E��K�۷�w�����r12�w{��E���r���J&cQ+#'hnȤu�(�[�jS���哓��Io�2,�%��SfK�'�86نĄ�= �9J�a"���>_;�v!��P���K
��O�|a�;��9��l���T����|�%�L8�C��ޤ��1<�"DgسD�T'�$�W��B��z���1���F�����ҎPx�4��/����'!���-r��-�����&���	� 4_<{�*0����ݥ�
�Z��(�|Vj �t�����Z,s�l�1��¡
e�Z���gM<��ߟ��$>b� �8(*�˓_�mHUq�ځ�J2����5��u���T��ng1�Ax�j33����fف�~R�l�x�<70!��z'�5U�ͧY!�T(�T-o���I:i��Q.��g%j/^=��
��K�)��r-6l�B���GU�ϸ85������*���:)Ѹ1`w�6$�Ѻ~���x�Z[?��ʈ���y �����k��s��UG�~��f����F0�a��s7��*8�#\I4��[V'�W�B���BP��qFK���46ӳ��ӗI��v9@�F��Q�K�o��W���&O���B
v6 <�eQ�����~��0_�7�d~�9���]�Ĵ�U�Ѧ��w��}K�������k��2)�^��.!Nz2*	���*&�rl��!�)؟`��B{�#�}PG�8�ݔ�z��e���CRc���}q=U�}�9�)�����6�	��w-�:OV���������l|s�	�|)#t</���k'a�K��f�-DeS44
ٙz�3�L{�<�xn�y�-������"�����h'���������t܄�.j�Jh��[o`~Y9n�T*!+�Gd��8B83`l#�`���l�{���a��o؅'u�5�w�>��Z������5�;M�5*Ю�=�L�3Ԃ�������t���+�=���?�F����%�Wn�8QϢ{���s|�A5�FnI;Iҗ!�����Vn�49F/����X�b*Z��|K����~�N�@S��[靟�~���i_؂�G䧖��`�� �Bu������~�^y�mfT㗈3Q�� �����s��>���AH�a�ǫ-�K�i�n����5�Y�tIzq�0���mt/_�S�T���7�W��I�� �X�t���<(1IDԝ�dZn�߅$5�V��S�^m�!V}�3��o4M��~\��k�p�˿-]�����=�r�$��" ���_JW
p�)G@�3�$�AA�ڂ9���BCbO�t����T.t�{�Z��"����z�P�Icz�Px�ai�}8���^A�ᅺ��N���q�E@����z�х
�@�WooYe�$��$�xD�nߴ\���FZ�d���KVYn��-b$���=HS�iS�n����,����|��	��hKi��d���fX��9�ͥ���x�^%��:��!E�M~��������sx] 2pX~3}��-'8L᝻$U�RuUOuU�9�i�S�ɾ;W��Ia���c�U}˝o�#��]#g��N�W�Xg�ˊhVMv��$R-�]	9w�������] P�^�ɖ��v�9�*͛%���x�砻|d5�k	��v�����ߥ(��3�<:��r�|��_yyS��/�KA"�O����6������f9�fR��n�$ͯb1j\��@��g"sQ�Y�j:Z�Z
a�Ӡ[r����hf�8�6�"�a��|7��K��c�o{�d���s���g۶|N�	�^$PJ�%k-l�NB�� �a�EY÷�1���+a����+ulGɻ���n�}H:���� �I�A�0���W�-4� w�T(qx	T�~cI�Z��j��UCvu|�1�p��셝	Jdꫲ%�4Y��l�}���U��F٤-��|k����ę|�k^9��Qվ��=�g����caX���];��L�:�0��07
<n!�W�Rr{��Oԛ�
�9����J*���N����
��hD��y
��a���qӠ�B�h���N�����؀�����.�"�f����(�~%�FN-*�����������oMB��UH�q/]�?U�n^S���CU:ۇ�V�;��=B�dUXEf��T�"EZg'�nz�N/1��p��0�U�E\�tS��x�����%j����=�W�ɡ���]��)��iܭ�f��d2��8i�Os��D�E�a6�}���u�U2��BS����n&N�6���[�=o��*v�,?:ό��;s�[�2`�F4��l����A��h�t���9r�bS�p�&^s��U�2/��ԌЄ���_R&G�����K����S�xʉ���>�Z�)P]'h����kP��� R�/�BNY�N�W���'-K�M�hb�����h�/i���+�Ԍ?x�� �2�2)��"Z��>���a:���Vj�����&��oSh;W[.���Δ�v�y���.r�͓�sZ��޷W�»�{^�p	r~r�:7�M���.鏱����J2G���Qg<�k��X�fNXv�KJ� N&��y>|5��
t,d� �<s��"��:�Srx�<��t}>5YBB�4X�5Ys����]��C)X���B�;. ���,mǕf�l���"� ��\`&z_]m~�I�P�s�	�f\�P�t��z
����E���xnWH���d��#�����e��*1!o���u+�}"��U/cB�ɣ,2�B��>���5�a��}39�����X�f���ܨ�(��w�OI��3�����Gd�Y���~��!�F���*����BĽ�_ߝ�8��3������G��O�?�F��f��y�6$ ��qvh
�f.��e�B��tab�܂f�UP���ha�g��!q�/���Rw[�@e�w����a}z��q��I7��r���)�DG��f��f��VAWC9>����\�	�죇��g�1᳁�y�[>����:;�E\��u�V���EX�D*�i�"7F�w�y���#��Lvh�銽��NI�z��)ߝxu�]��F��U&U�mcZ/����J�_R"�F��Di��u�*��������˂���9:{�u�~��R��t����=���Ȫ0�{���",�!k��'�܁��4:6[�7�6S���2��'hm��3�^������ޱ�Go�Aċ/ƞ�c��9�`9�*a�y�L��6F?� <�[£�N^�LW`�[l��i��V���\������}S�����%O2%�J��Da��}��OX��^�a",�Gr�Y����.�%�	ǈ#݀�q�?��lNZtYlRH(�oa��Q��&��D)Q4�Ќjggpj=ŋ��w�T���ٙ�Ĕ�}������\�e�v�g���L����"غ�HFV-o�P�e�8=,��}������8���ҋ�ޛ8%t�ړ��.�~�����v������=�_�)����^��f2F��/O	��ge��V����t�%�v�F�I�8��EJ翪eD�$E��Qε������F�^�!�W��bXH�n�?ɹۛ|PФ|�N3S'�1�:^mB�]��D������Kw��+�_R����U9�f�(��џ-�u��K��BC��i�'���������e���59+M?�LxS�
I��%�ُ	����H��ݵ���	��R�K�i�@~r4�Ƈ �ۊu�����^V���'ޢe�>��������P|�B>ȟ8��x���y��ni�{�,��	Y�:ʢ���H�kFr�VG�Z�\}�4ת52�$������9��E�MM;Q���#��>Q:��\4��Cq4��ɗ|���\��,�m�3@�g���La����7�{��h�l��Ğ��M�(l��/�(/Z:-�k� S�MFLsz�_��"n�+�~��iA�H��^�!
X
V��h�%KI)�(����{m��3䝧Z����C���M뜄���(2P_H�������$�x�L������1��!�5;9��&
吨o<X�:J��Z��� ���:"_��Tvv�9g	��I��>�ٝ/���B��g^s{�k�^J���	�c�鞛�q�d10��L��
�>)?)}y�4���l7���97���4���O��"��jt���p9J$�yS�YW�,Z��E)�v��ZD�����4>���s8i&Gj�UЂQ��i���7��v<��D��
9��YU�U¹8��C;�V���.�l��x��9I�N�5���x��L���a�K[	�g���ӵ-[�\�؉^e&r�7�:��dj�>�$�k�9��u��P[�*���L�w��	�w6��}�֟. ro*���F�;R����틆�~�tf�)��Is�����Xs�9���� j�mZb���}��}��́F�%��E�7�AZ^��_�w�@�P~Yc�c��"��x-�W�L��⟃���P\Oy��QcN�1_�1Ꭻ�!_ɐ�e\Pȍ���Y�������J�L�eB>d��З�Y��<'���Q��R�E���RCx�ʘ^��φ;���믦6�g��4Nպw������e���೸��|pP�8M^���4B����?�/P�A|�Z����4{_�JᎽ��U9�:(���Zv���(�o�<(���h"p; ��	pԯ����Q�B��7�gLx/�l�Q�Q�9_+A�?��}C�8��/��XwśR�"��� ���a��Ϛc.J9�>/����Q(�"���!&}wAv����;$��m��YA���1;�����6��p�='e��	D�.S�x2�e�1�滣r�sLô7��[2�e��~ma0��m':# ��t7�r���%�n|�g%�ӛ�+RͼAР@��UϚ�ǌ���T_K����ltL��|�,��<���<�#���/TS�1R�Wf����k�E�\�P=�9٨�;K��^��hp���������a'EЈ�A��;0���ef�M�}��b����$�i��u����yf7{dܿa���R�_MIZQ���^�k�Q��,@����oXk���۝Z>��W�y|�qz'-����QE@�`8@�"w��X��D*h�s1�^}�aL�'�#�<m�o���&�-�F�.�&e��8^�B�T=g�;8��F�=ޔA;�S��,B$)�u�}�%�g'WN���M��ٗt�ܡ���D�M֟���V��j�׵�&owyb�V\&Xu�T������iGe����cɅPXO���f�^�	��M�YZms���2�-R^Ұ@��F't?��X������mۑ}ό-`$)@I����ԝS���M��7��ޛ$�(fm� ��u���=�y�8�} #]@r�%���`x�`%PeNV/�'O ���sOƴn-y��\�I�r��P�i~�aW̲Ȉ���L*W�ќ}�ʬ������FԸ�C�Kɮ��8'kMc�3�/��XWg"�j�r^��5c��q�gX��qU-7� ���"T��,|����*�^��Sy@���k�'�u<q����)l�>�q1�&Q�������b=����>��I�,b8����|�fx�\��ɽ�gO�<�
C�N���ǽ^G1���צ�OP;Hl�A�ǥv����ƻ�h5�h��E�2���
ϸ�Ҟ��f�v���) �x�ʹ]��wx�P)7��:r�5֋�����j��pz2�2�\RN��v4n�%{��>��>n��O�j�͜W�5ڽ�Y�n�M��������	%��h�T٬���E�sŮ�p�"�r0�[�u�7kɻ�r>���wCT+Ww�;S�[��D�zX���	;�����s8浹ö�ɠ_�˳������O	��w��.�~��s��2�9���H����x!z�)6�l4HY�I�#�7�PK   �M�Z?��O�o  �o  /   images/ffe61187-e64a-4024-8cee-95dd034d2257.png -@ҿ�PNG

   IHDR   d   �   ��z   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  opIDATx��}`���ݽ&�ԛe˽�;lӻ�5���P�$$��z�!�)�1��ƽɲlKV�~����۽��tw�-������v�yS߼y��:���?����V���O�q�J=~��g
~F��1:8l�p�	�1�A~.��"8�� ��W��b�l���@���s3h������az?zz� �S�?���r��=�|��@e=֑#��!� 7/��j�����3���7�,zz�-���	�+pЫ��p���Ҥ�~�c�͢�ഡ���g�dE��I�7�~?�=���
�dQ���i�9�XY��o����&g���QD&@~푱���(�`�$&�.��긌�O%4<����ϴ���2]���/��h���0�=�Ֆ�ȴl�}=CI�cJ�3��6�	+������ޫ+����~W����YPS�"6�5�pwց�*�F��S��t��e|���VI ����XY|^�������g�}hh��>��|,�
��}0 IAB�P�$BN�vR�JP�]P��Q��>K*`�M`
-Ha��Gp�"r�2ɪ�}3�p�7�O�A��{�;.��,��(2km䢸`���b�	���Q" �o���Or�@�ߤ����z>�i�g��B}36�"!\��@��U#-T�15��%�CH��N��&�q4�wkJ����~s�#1���§W5¨,�M���@�f㳼��e^8�7\�0lLU��5�T���F8g���V����E�L��ϧ�a�����SjC,�ק���1VUd�&�{��	ɦ*�M*{^|N�>���=5.�}��T��Ќ�B�.���VH����7@�dO�P�n5�]�Y���9cݰPl�s�I�N�^	�y��3d�� ����ۀU&���<��� f��ŵb���\����b�"_�T�}���p�>A��gnY~ %&+��=���³V��ML|Ρ��}�GU�c��j%�=|T6�BiU)>�ϝc���-�@�;�ꏽ($QPg�)�7�>�^��Qn�g��Z�o����\p�;�6��(�� }�k~����� *��2�e��������Z�ʄØ+	�����g���{��E��c�2�c*��)�-W��A�}p�0�2HC�7@�/��&���f:T�>H,��Ud���c�
<6���}�^�d�FG/d�	����W$�~|�����Zdܺ*}i}�Ow�p|��/&\�����[���D5̝��������lcO��x�Y�>ϭ*wa���h#�q�@�e��<>��Y#��$*��[�����'�破Q�X<��2TRˑk��
�[�HV`j�~�5A��Ӳ=�G�z� h���ށ��;�f|��	2�6ݩ���u" �pq�l)4��! ��OH}Ы�{q��ע)3��H½���Y~P�gB"9.d���^D���4a��Q��u���U%PPsI)��a������AZ�(�I���EC 9F%��ټ�E�g$ꞟ��zGX1pS�8Be�^e8���w#{�!�l�a�7^��D���a��� \�%�J7�w�]�$c�_m�Fl�����ή2	����>w\i}5���'�Ҹg�܀>B�ۡ�c>��d7ͭM�&b�F1@�O��ᶩN4�;Ψ:��-m��V@�(pKN�����
�K{?��F�	B����27�B�lwGO��r�A�������&:�������bl�%C2=[m݄�g��'�ɲ���@vU$�Pw�N3M�U4��F~��$��Qj�CjV?~�'�h�&�/w��MBX+KDMi4���ê5(� #F�뮹|(*e��#�R�$���s��;���9�g�Yg�����~L/5�;+ެ�E=Q�).�O?\��hdX�o����_^i�����h����L����a_���)��K�n���ݑsF�/E�/lB��S;h�7��T�;p>*����o;"i�mP��+*�j���B��|عs/2"�8x�b,fHMM�:�[�&ޯ��������?*Z��0|�`N�����a���J��>En���N��6�U��0�G{���<�ѻ�/_W��Cv( {���wyF(A���� )k���dp%'ˋe����jQ����n�'$Ҋ<�TH�����RB���_��u�Lbl��*(�?���|d����Ñ��Px����W�����X������U�a���p�ݷ���'�ۊCF8�&@�	���*s���'���4����Em��^����:��Ҽ�V�A�`�­�֡�V.���Y������K��)\�%����kVc�-��<��o6^>�w�q�x��8-����$''�����M��$Z��=�E��y�^M�5t�4��H\ѳ�+�����Oq0g��sI5D���W�wz7�b��@��#�c9N"�W�8[S� �D&�cU��CB��P�Wz\ቂ�����&�=�ڹCE�'g	��n*JZ��EV�Fl��^�.��<HII�%K~��*��\�������l>]�5���~p�/Eb����s-�8A�P}2���N�S�i
��b_��8��
�\��;,���V�%h�]o�o�F3ģ���?�X��E��2F0>�ǫ*F4{��2@;�l"R���_��o㠰G�<�&�ڈ�3��f��,��d�F�4�l���#�N�1��b��Ǖ�r����l<[������0W���C�9hP8���8����k���A.:�<$z}���Dp5*���m��}t��w���j�#�����&QE����hxB���+S�`rl}G�þP$��N��;��I�GUP�A�x�����l�/cQ]L:͐WQ�GG��/���E{�p�8�A�O<:V����"|�r�k$��.D FP�D"+>�
7\G�ǟ~&$Tn�����⪶��#8TlQ4��=���87T�H�K.>���p���g��A	���D����n8k���H&py��
�p��)0{�P�);�M�����ol.���	���a�K�o����u>����U���<D�k�WUoC�����Xm��mHe?�>UpbL��?7�C��獛	ŵ��5Qƴ�����?
�`j	���&M8z,�"�qDY���e"��'Z� �VyME-�K��MLM��@;�*�=R��=QA�e���M?�,�^6��>�l��XZ����s)�"2�A��sƞ���?�qО9�$�j�r@���q�$5'
;e��:�D�I�d!9�tq`��U���r���D3���K�Ez%X~�]8�,���]��ӝMI�������x���� ��MK�M�ε ����½P�WFNqCg�D�煿@��F
���o�&?>�Z�4KJ�N�4Ձ�h'�FI28�/Ě,��#H8�$9�1ML:����&v"�dW�D+aA1z�B"�\�R�ϐj����\���b���_	K���x5�H�A@ܠ2�a�Ep���Pଆ)	bM�Y��|l����$�� r���@��?]�1S720(��?��5�s��i{�������i��}�=��Ͽo?���I>:����?��&�i��2$����%�����R1��	�6%|`��M�q6�P<ƍ�ښ�t��d����O��专�_�_@��J�H!DBD4d(m�uL Hڧ+�v"��d����=��^wh'�S|YW)�a�ps�f� V�UBo���־���J�'���A�4�N��~���bI�^�!XYm:G-^�np+�����E� ��&�G��,Q�4�e�dM>/<_Q#�q1ɒa@ب�1f�K;e����nuX��,��#�0��0'��`�bH����&�E��
���u��(0���h��c�Ǘ���	>��򬲁d�ǲ:�/���5�Ϛϐ�D�+v�{�Wv5�~������!;�C�֭ �,pY(߁����,����`��<d{�.�!�s+�B�dUg�`B�o�_�$N=c�[Pz���A%�A`a�E��Ų:p�p�D��!�aGI�2R3��q���-w��S����H>l:���L��	:��0؎��4hlD%������tn��.��N��&g�,͇�Ź�x^�#
�#�U5H��lF�*�\�:_��h�����#`_y��GɌO���x(#��5,=�[sGL��yy}uk���@�%��	��a���p"�ݸ������+�y������G����	���t�QĐ�J"F��&]b0���t�F=��Qn�=t�I>��g���Z�4��[���{�&�C")5���˺��"to��� �>��{�WM=���xrВb��	O���ѳ��蠜,~�9Pd+�e����s�Hx��[�
^�?o�g"R�1Brq��火���n]�mr�}Ӡ��:Lv����J(�)�8b�YӠ�����	�)i)P-�x���0Mh~S��qEzdp� 蓀m���6�hn��%@Ecm��P߲�)P[Yퟦ��48�����T�p܎��w��A�?��O+=��[��Ы�k��^��Eވ���'�?M�w6|�G)!����/�DF3,ݻ��hq{�QC7�9���)4;������χ��۠��+�u��O�������Q�ז��h��Q\��_�X��h �;��б�6x|��;��p ��?ݷ�G��#�U����$�Sƻ�|�I����&N���S�(2�q2� @QeQ^]D�k�E} ����	�W��2ma���nW��	�G�n�'�~?�Ǳs����<џ�7��O�B3)2��N	�5A�qb_j|�.R��c&�gA�)z,���&�R�+[��>.8e�'�(%�#��Q�M^��#4�@��_�z��S"pU����t��t���A�D�������N�3�_�8xV�7YJ�=�s�ֱ�d���w4�?,�5�r�1r�[}�����	e\$:�9��ף�36.
Q��q�4y�Y��	I�+����/C����H�;�k�����D�	*��&I�����=���*F������v��^��j��R00�������n��<��pEl3)!NA��F�;њs���ʒ�/���p.��Ɨ�C\�\v�Y�c'�>�%�+)s3�;Y��gE���î�"FWھ?��,��cgK*q�r�'#O����������F�W�k���
��.a�Z<���;$�Q�Jf�WEٽ*�h�]d��^�>p,<2�rش�4�|������9W�}?�;Kr[���dr-
54Ei玉�O/�{ecu�}$���wa,��N�mMu�:��Ip�Q���_��o�a�*��/ �?&��z3T���?��t�Ȳ�S�Z�r����ϛiB�/@Ѹ(��h�#� te,+(��AY!|.��Kђc;"��נ���׆�߹�R�{��t��#+�8X��c�YjS��׌��9���:��5.�G���y�0��}��1B8<�s�(����҈�C�_8p�;Cen��fZ�k��&�n��*u�fԣ�-L�V�8�rZ�\KI��j�����ֽC��8Ś���j_�!�^�J���63��GH��b$q��ə�@����G~�>���"��zb: �ÿ����x��f(�v��xTB��>�� P:�Q���;��楂ݨ��Jl;Ú��M5\iw�H�PTl)���4qNo������'��&ua"������O�1�4����W�R�{$��z3��Zc{$��;UByC����_�Z�^�!R��HKi���a�8}Ѽg��isS�O�=�;�����\�fw���+5c!\w�F��,chىh3��Ɵ$��+���#��V��N�9Yt3рh!�k��R��� bг���Y�qM��M���[K<.�'m�BZ:���>�`D� >2��H�[V�Mլ��	Q!�]gE$^W���V����7W}И&�#A���T!��צE�5 �8�m9�pF�K7�nm�}?�U�T�Y"k��0Ev���V��;P�Oy�xl�=~�'I�eW6�E+�@�kp��� 5�<�?��"q�~�/�p��LY�8���a�y��!^ji�!����>q����D!�T�P-Cz��Hד�¾=y�1���;�.�`��e4�ğ�A��gZk����M��K��oM�(<i�U�( pJ��[�<r=��$QeCu �Ac��\�W8��i�{jjj���D�L���Q!.6���H)�~���6bq��E���\,|�#�!��ґ�F�^F��j*p`���L�M�N��J����!�|�U>��G�?Z,�u@t�?{�,(���ꗘ��w��&����
Y	��i�O3���������<n���s�����Cae+Az�l'r���(�qDuW�eQ��N<���f�~޿E?��Wь���Zp��0b��V+��1 )%���������Z]��.�eI�|�2XlX��߇�Qt�x���8Y�� dG���DN("J����l�R���@�VE豬H���+F{��� ����{K��,)-��q�h�V+477C^^^��s��U4-���a����F=������?ڣ�;k�IPX[c�PLaM���lHg��&���u�_C
B6�$3w:�?�i����3�����B�dG%���V7ќ|t+kr�̡ཌྷ��$
���%d1���@G�������>��l4h�X�!�}��v0�D33v3c��h�����w�DäkR�R>�q5e#F�A����r�r��-#^����so�/����I�j�@R*�3hLmST�z|�s������O��p)�.� ���;��]�u_�n0�$&|��0ۚ� E}#Nɢ"�h�|�)/���\}���x�RRt�f������x��F����������zgL�X�>���&A�,y����~� Uop0�`�-o�����d�7O���)����lE�"�u��>�t�zm�pO����d�}��B�+K,��D%�qg�;�D��Mu0/>ŇX<:A�DJV�2�᪖}��^`�GUO�������6�5�o(���dUD����o�:@i?$��EVO���T�S�6=��RA�{���	�f�ϩ��XO�m@8#ܥ�7Tz���.���(16'p=��~]_��eɦ�+caV���ld���Z$ưZ�w��m~�,/ k\X�P��6��hK�v	)U�
a��תD$�~� 3TGsj;�/8v����e!���vl�/
�Lټ����|ދ��7���J[7$	��|�e�G]P�_�	�e&��M 7^C��g[n��GS�,���>Z�#2���N�C�(F��U[��W���ZE�ar��U�b����͋�J���HEJ��[�#������K!r�,�yG31{8��n1���w�_�+49��9b.��	q�����z:�Z$����q�i��,�Ӻp3�9�)fO<�꒮�\��]��P�0|mVu�^V(�(9 ��\�����C���-������BjzZ�*>�@�F��s���|"'���
�����́�hi@���jeti,e�}��������FmC_����				PYYɿG
�P�dРA`Z�+](z� tQ��ZH��B3�59�}��>əPUUŉ����z�����п^d��-��� *��2��D�$��P�O:�<7�-�x���ƗF���CEy�; i(���%P���zp����^qL���o��C#�2�%
Z,��g�^f�5��kFD�Dv���]����lXͨ�o>�T�q\�qr�$��|�!�u�PU_ó��$�Y�x�7>S@ԇ�Q!_�y��L�d䎚,�Ů�@�.h�H3�$�tN����fbY}T�����w`G��4X������4i�9�&����9:Q�>)u�9��7�������!Ȱ&��P7����q��[�-ű(���v:[p �]XW�m�
*Ø�*_����;�*�Ѕ\��9ݚ7�e�;���,-'kfp34&��F����NEYo��g:#z��e��XQ��E`��	i��lk���)���~ˢ�N����D"�\v��&p�+�Ԗv]a~�=�Ó�K��#�]U��<9qG8|Y���ͮ��
�V|;��B�,��jɥŲȃ�eڶG{�H�x5�����:� �/�E�Úo��Q}��~Z�W���W&	��"o�~Q8�^I�j�N3תŲ֑>N�4���%{A'�h@sOR6�)� b��Q�aM�7���_��^���*��m<� @1u��i����}�"g��|K��g�h�ꄻT��ʛ������M��j���)-� ?��$��.���,H�#d[�l��ۯ�s*�i��W�kmŚ�g�@�����@������p��h���߼�M�����L�3�h��벪^ *�E�(^����*�A_$��H�5�uPJK���~4S�\	�8��i_)W{����A��9R�3*T}a��y���N<�V�Lk�d�0��1��bF�z�|��׭�VkyY��e1p�]�t9[^���C �n:�B�ڗ��d�d���z��a ��x���3`|�`ȩ9���m��x�Oܔ�	��CA��@����I��ՠ�܁��cP����Tmo��6~�	$)C�)Lh�P��
V�W�>�����Bx?�#�,��ƒ�~@K���>o���d�WR�6��b!"��8z����êO���
�A�� �͝��S,Z&uW�PP�jk��Y/kӱ4ge@�M��6�^qj�� S�|Jն���B[{h�!"�o��NZ'��a��O�Ao������9B��Y�p��&kV$c��)0ޔ��*��F�z��i�X�t���\���W ����Z�G;A��'_I�X��ʏy ~��F�RSz�i������:8'C��I�,0����c�an|J��5�����ʄg��r=�3	i����x|�(K�%oT�T������Ñ� �	�(�k}���"a�8r��_`�޵�0KQu)U�����N�M�ߥ�� |�?w��~)���DK�L�.%���T��&A�.p�����c�*�7�LL�q'rIg�$�$�^��Ce�<�VD4n*&��s���(���-|ݛ(T��}�r��w���1�ť���k���A��$����x�E�F*W父�-*�Д�Yj�v蕀��֛R�W���z��\�hrۏ��Ҷ]M��iP�d03��ZE�,7XkUH�5vTR�HH�O�eMs�J6,K��}5��3-K�]�\���@��'=�9��53�����ǧ T����Z,�p�b0^�,��͞=�[��ZZA:�9#N�����o�ȿ<=�&R,k�K��!�����%:<ͫ��d�Ɍ,/�����?��Hj�[pI�S>r�}߾ڪ
�?t�Q^��
n3�o���f���x��"�����3�rU���v������F}���(� kNIfM�
W#�x�G^�&%"©ԑ=Q�#Í=�)���#��"�P������3P|��/iu/t���'�$}�u�9E�<~��c�C"�ߵ��l���M����*_b� nKg�w�=�{����1m�I:��yYv-�xQRD�to��B+��w�e9Ƕ�� ��{�lWڼ��f{��6ӱ#xd�}�,A�4���	�S�	^(˷N���s.u��@e��1p��S��� /�,��Ei�� ���?�	��H��B��'H��Y���A~B�{CM>l�/�y��c�]z'4fD	"�͂o�Bz��C\`0�32�Y���s��k1�!R߯)W�)*��[Y����Q$RRb�u�� N��T!lUR����2�=f����,	itU�x�X�ɼFth�H�H���qԠr�7�B�h 2,G\�A�t��oEX"��Y�Id�z�"/51aa�m�ԫ*sЉ)��M�?���G��&"
-��_L����O�D�*�����z�%��mܪ�[�(}&5Se߇Ĳ6"�J)�\}���u� H�Q(�e��z��i������/ ��"¥�q9S��_B�����FtJ%��ԙ�:ѩ(Ih���\XN;���tgI�r�"z ��k�����8D\~�G{�L�p���kaF� �H��f&�6D��Dq�r!ʻQ�]!�>@"WUW�ּ���A��/����v�c�h۾N�O�nF�Dفz�r�!t3��mޖ�T����Ak����s��q����`dЬ�H+!;	�@��R��!9��������Q>�8�HY7Wi<<T?b:���o���	DI�V%o�_?�8Ύx\�$��W��	gզ�(z@Z�u�T�M���
�m����>}औL�gn(�-�(V%(���9t���D\vJϤ��n2 Gg�j[=ז���!<����%X�`d� ȯ*��Gg_�7~n�w��$�����u��Ⱥ/�E���$��u$�b�ŭ?���90{�$8��D(���K����F��XT�֗�[<Ӊ�E�Y;p3\cתQu%� Jg o��0A]V
�I=ȸ�`�cR�Hi�ym�������[�����Ǟߕ����'�m��!����M0�2�Z8,Ԁ�t��g�����J0���Y��/JCi��,�� `4@������pZ�KƉ<Qc�_�Ѯ@�P�&z��I�Y��!ǰ7]�t��U�C�-f/�ߞ���}�{�W�@����7->���xE�5kւ���9�p��>ْUc��22	<診���.�h�����0Y0�$NKN��x�阗��hթy"���I�]�$�'�En��X*�JLL�~������#�_�Q�((/��c�B�lB� RS`��q��Tղ��I!�n���7(o�^JC�A/�Fb/����Sx4BU�>�<6%ů�lN��\�r{�0Xok���r���i���57�s��I�����[��g���E��L+��XW�~�2b:T֖�Z�ڈAbHF�6	u�����;i�}�x(u��K�?�ha�5�B��
_�o��5y����f�p^������ږ��bY���k�렬����(�H!�DE�/�����4+
����m��B��6T���^�R�޶j!';%,L�����p.O�얍�X�r��ؖ�rm��(aSs!��Vr�A��2�U����lv�� ��L�~�$-�����,�4D�e��g`GCs�+�˰#��%N~����!
�|~�����L8�/�u^.�d����#�7����]h��(�=D��Vm�V�����ے�Z��/?E�`�!�X�#c m.��GLц`��#�<,��(��r~�⻑r�ZNB�OU��{��0Û}uAR�Ϻ
�>G�GK��Hɑ�v�� a�	D!iۑ�7�qG�X�Ze�E7�e�U!1�F�6��Q�ۓ%�[R"����xP�d-#ٚn���(C2^���8��Sa���P�TFd�ԸDx����2x5k�l�0	׽@r�r��Ғ qG�ŏ�K�N+��<䒵��b�����������H*5�JzB�쳠A� � lF3��6�_�S�L�g�}e�� �o9�:�o(�L�P��@���A���� Q֘�o���;�ċ��C��@����#�q���8q�y"ݎ���ZZ��m0�"�k	#D��{���1��� ���� �1	��-�q��m��������Й��%�����{�RM�"7%��<���j^�!9!ds|����8��&Z�3�BU���"�0f�Z@�ά#��nH�w�҈~�6I2\�o:*��h�#���dS���ǡ��C��ʦ�2���!l)ʁD45�>���3zee_�Z4��A�dn�c�C^�=�&<9���
Vs`�V���P�:ѧ�&���h��k!��z{���a��Ŀ�O�.5��bY�k�S>j��S�(>�j��6��^\W/Ք���8Mj]˝̞�%��AN�z�<�+�PS[
Yæ�6~�5��n� ^h@o�5�7�ldK�:@�`oh�)�?�ᆑ_F��T�m��q�HJ�!
�����*�[S ���:�d��![=8z�o��R�{�ύ��5�Gx��N[�{�#�$Р��Z,+j�\4��t���a���Є>�+�I����~�s7�p��S�Jk���À����~�=%��t{�.4Kr���qr8_�z�8L�0�d3�䘬�����!�h��g_��/�i�
Б�SQb���k!=d
��K�8%_rֲә�
���I�|$�%���B4wq�k0���q�`���6-���7]y`;��%@ay!<���S�����j��w[I.l����-�F�N��p���!�[vt���$��#�?f$I"~$^}�ǡ��:>��N3���~m���jQaoDT�*���b��q�p��Oj��Ъ;�
�X��0Ā񂨥��j'������,Y�����H1az\��զ��e�+&��@-H�k��a���/xp�Lk��W�+q;���%�ǲ�	d���q	�d;q�_T�.��4�(����a�@bd�b���TL� �� :�$�j�-��EJ���}��ы|.�|=������9$&�`Z|Qr��i�)�a4�<���|�"�em*���wah�{��&x�/!^�	B@=�N��Ę���0⎈���� 9ā��d��� ���GU�l�{^*B�������fz�q|��Fƶ��:�d�*��2��k�� 	�[f_�'^���[g-�7�-��##��h��(��[�vt��嗾�1:s]�3�Ųތ%���0S�V��J��j�ݭ�����f�h/x@�Z�АB�SDb�(H����zO��Y�i�����+�Q}r%�]�L���\nXbL�@>�_��8Fp:ܜPԖ8�KA�1�W� �3�]
�#.2Y����b�SI�3%�6��#QD����_
��C�,l|�jt��촃�__�\ҹpŤ�|:uKQ.�;���'�@�N:ÇD�XL\d:bb����8�d6p}C���AXp�{��S�g��3n�?��g��kR��+2�c ld��uv�:u4����~O����~��
-L��D��ZXE���(tJk�់_�,+U��u����P4��C<��'� ��8�5� 11������>�lX��b��\|>����'��p��"�_�8#��������D�e!�@��-}�q�<o)L�w:@�捶O@�G�[�����T\���!��;�9T��g�l���-&�^�kDh��
&h<0�ɆX0�{�G��5|*���Q�X�o����E*w}z�l4�I�'��R4��g� ��	eu�]n`LdC�E�)K�����ne����22Y�o���(̐�f.�U�oc��@I�r!Jc��ѫE-`�ʺu�\�����ҽ�!3!�ω�uQ�@����!���"�n�:1j��脢�ta��e� 2Qg1͂��p@���w�$i��z��R�A�%^\�Mp��+`����ܲO�ˁ��("H\9Њ"L�m���r����p�BD"�ߥa���~�h�����G��}�Jhvt����ˊV�'R2 M�o][6^Z�	��[�T���Q�YQ4�)hH[b�@���(�z��1����J�p�t�zq4;q  �/�9*�7B3�fbќa5�+��yY�$#;=I�*iP"~'Χ:[�`�[4*���zVc��W�+�v��N
�������oF.p3�]MF)PƜ�	�}u�?T�lW^ }�B����E�:_�}�C7`rl$�_ş��z�c1>�&��^��>&��\��4�=7>%�bY�WX�h�ѧ�3D0y�>c7c�Ez�r""��ڿL���������4����@M�l�^=�
�?_d��}�0�y,���\��(�Zx��$H�����.���E�c��6*�6�ٗ��hY|qr�Wå�#���}I�6��yy��Ě>hL1[�������s���ُ2�K�w�<\t�xLK���%�H\Lu����ט�δq�����τRڟMD��p}��{A�(ՠ+q*:���8���v��o?"=�q�̋*���mS�K,70a��Z�ƫ*��7ZfX��~�lcm����-@��������ִ�#���ΊK�2�a��Q����ƴ'ӱ��G(y�Ũ��*\�wm�[�͂��}	e���a��X@F'�?U�F��pj��2_�˝o�U-���y���i3P�� j!dMB���"$B�E��� b���x���6@bR:\5�t����)���(��n�_�׋Re)��N	b'���*D�{M�4�^w�/���c��'�����̈o��f[C���o�����#Qƃ��S��ޕ{Yk���~�:��ǎ���(G⨟�o:6��Ecu�xM�����D&�}A�K��t��8��9UO��+m��f����RF�Yl�Y�Q�p�Zp��������w���w�D!��.K�s?>�JdnC�ވo?%��	i���Gh���k�o�߸����?��o�<WK{� �O5����l��@Z�;�yH�G )k�ь��B�Z����uB�d��9���m������F����;�$W��v���U�`M*7��u�1p4>�pg`,�k�s��a�Ixx1_cx����e�f��ݎH#o�<o��^:��K�{oYTR��c�Q�{]���_�A$�9�E0����@h������-�v��c�>��,A����
b[r�1����	R��J�/�^��?�9���RT�F��E�J�J'&�����c>9 ^���H�u�|�&�d_k.��<o�Q����)ZҠ�����h�����X�� "@�4���hL�lg��I��*�O�\��i�;�s���\w��n M���^��>?.�s�V�+�':�_m����I�(��;�?C��ޞ����9��`,���a�Q�G.)m>��X ����u��Vŷ�Z�l}��ߙ�M���H����F�(�5U2�	im�R�e�q6�[���x�
p��O��e��,�4�K����i���mus�,(~�/�B����]�o�&t�Z"�e1zc"H����Br��anCS�yxa�B�#�b����ke�E���d}�q*���[[��uK�c-���M\��K&tw���l0­�`�)��Y��tm���
�R��;��(���{�ιdU�򶌁_�RY4h�9v���}&�QY���8�2��yW��%h�ъ*w$��@m��	B�-G )�1w�Vb4@��pg��[p[ڀ�׫�/D��&�F��<s�n���%�����+���[دeFA����B��_���l�y�M,�@��Ef���9ẹW�)C���:�yR��������p��#�?�8.|���r�����2�����]�R��1�.	QWkN���ݺ.͠�hr8%���@U	�?n&Kφ�YC`���G7A�_���U��8$\J����F��Z$�#�Dj%l{�A`�ă��'7˾�D-�u�Ą���@a;r��MPgo���WV����ˢ{ g���2D�V��@�E�����YPe�)+�_��"���w��Ef+m���C�x�;
��=g��ν�9@��,��<-.�}#�Q��͖̀��j��\��J7�4��_UAk�@�b /z�1&�ڏy��т�R���w-�ڛ�8^@bka������B�/m%��ɤ
4ދ��D4�<������'_ k�w@>rȩcO���P�uG:i+PU> �d��+�r���~�!������F��
�z��?O��fW%�Nw*����h��'͇��)0w�xo�w�|!�	2V�E�s$.��R���8����K8���.�e��C&�9cN���#��m�awI���#d!".�	5�\dUWBIsJ�.X9���R;`{��i��wۗk� 9n0����	�����"�҃��>�S��x� M��O�/I�OCGp�_c8N�X�59���@[�@���B��t--C�KH	L�c;�q�<�Ar�s�󠲹�+��hr��7C��w��N~ބ�$*F��.h�1�<�X+��Maa"Dx��MA=cn�� �iC�%���Π$����G�ʗW}%�e��0�3%�Y���q8eb{\��`b"\�:-�>��]أZ�]߶Q;�bM�R�"��e���tދs�SU>51aRw!��#�<_xю���*��=@H��z���[v�y(e.w�J�E�@C�?x���F}���yP�aB-��Fֺ����(/�(��(���]�����o�}!ħ2��mR/~EJ�p(�E�� 	@;�I��M�V�P+�{�Y�螙�c-/�1*O(�>|"��z8D��n���A����I*��?n�g� �!�T�֊b�L�FN�f��F#w<A�r�`�KQ���:NUكa�N�53/��5h�ȋ+?���C]��������}��~B�$AJB"�x�\x}��=�� �������Y�t:N��WQ�̌�d�⤭����C@���8m �O��J|R��0w�d�Xǁ�z�YY�&��!�g��I]��A˥c�4�<��}$U��6䭚C��m�5�b�[*���cY-��`f���R�����rz�8�*=9M�!i}ᥕ�w���BYC,C3�vD�?wX|�.�q\������U� ��v�m,_[�.I*Vdu�˦/hߵo��^�U�6��,�Ԭ�=O�xϫU/���J;�
,���.�@���cm�%D��-x�@�W��?D���'!�~t������B�e���xQD�Kʀ?Ͻb���H���x8^�e�sf|
�m楰�� ޤ��y�2b�,=�B��a��̱	-��[���a/���1�u�ׇ��
H�����cf��"���>�����ᲃ��Z��?��jri�h��D^�=Yз`)f�ΖL!�L�;5�RJ��hf�֔�3̎��q�|���?�)���P�[��p�:��FnR���'�5�[�D4�Q�]����XU� ��|bؖ���l�2ڨ�'�9�,����dUy����S��GN�I͑��
3�N�kBN5�#����Y�k��'>�5*p�����	 e���>��x!�f�a�C����>��uhH=A����gNY~ �,V�S�{D&��g��=��{Ρ�N�xT��11�W)�U�S�y�K��a�A��,���O�����o O����p����'	��11�9���ʹ]+�H�{L�P����6�A�Q���<�B&)��`�d���iQ�n�K��)9�w�}��A�^6�S�y�O/��&-��`�[U������F&<�㰵M���H��#�@yS-�P�p�e�������[����K�B�%�p7?!�A�*�E��C�^�"k^P�x	��NE~P�2!����&��؋����/���� ~E���7*��N>�d�z�����_�Ob�u�E �VB�v`�z��Tz���
��$�%J��1���F�5��n����ūPd�/}�sǕ�Ws�7AH��DzU#'��bCR��;����#`���P�h������l�y_(O���J1*�l��ʋ�Ж�Q%���1Q2$��t�&w��'��~�
(L�@�(�gr+�xEk����z�̻^]MS�AV�����@�����e��M�/��;��6t�px�^7����ᮀ�jDvU��ǲ�ر<G��������B�,���x~r�6��/i���}���#��_c�$���C�Ĳ�
1��*[�k��p�у���AD����!�X�ǲ�"S̱�� ��	Mְe����2M��e%H ]h0),c�Ж;�>�xUŸ��ז�t����'��+J:��U�Y0)6�������[���RՉ������rE��m���ώOyݦ�_Ҵl(� �)��X������Nsga��L�o+�:���%_��s�K�3v���=�O� �a�K�o��.t'~���_��ɪ��WQ����p��&0q/�SU��-���L�>ź������mˍ#��'g��SN��J�P���M[�r"�/�cL<O��~�+Bs��T6T����z��oB*_�e����>E8�r*��C5}'�n$�����2M�c����NE��O�ͻ`���m���$�Ped ��TcV[O���z�D[3���`#�~{�y��Ew@.��w{~��w��x�:�"�©g��*i�b�5	b���
�3��;Uᦝߞ[�	,ܶ|nW�؟y�O��.���>����L��+Oy�7�BaM_���.���!���ֲ�3v�<��y5��j楬X���M�c���($�ϵEYh�0� ����p�	'���x*�k�+��w���|J;"	��Ms.���^'d���|��G���AA�H����0 %������]p\�������|�g�h��w���C����6��=�`g��-/#"�Wډt��SyA�/�:�:xc�bx�珺ŷ!��fYS��V|��3H�.G"��w����!)U��CPF����#i9�fˢ���OD ��?�TZ�$j{��Zu�#�,$g�#F�W��W�)g��z�z�rD���v��[�~(ή�r���`�swp]t��I����^r���c�jT!������"�Q��|�F�n�]�d5���"�(o�M��[-�i�ϓ^�"@�e�FJ��T&�҄|��VN�O���������IK*y��a2C�3Y���N+���j��&��\�*$!����`=��i�N�1�\�E����1���$��КuUi���gH\���^�������W�Hs�%Y2�k���i�']�)��<�� �ƒ�XV�����B�Q������3�JQ2�,��!�HE��>��g��5���qk�hi�#���Ӈ��W���s���-�0�^����
3FNF}d���gU�"1�y��Ho�)w� �u4A�(*��*,�.����Ew�D����������@���4��S�5$pYV��h�U�٣g���KQ7,߻>�m_�Pq���;u�/-���]2�,���^����Z�D^k�V�&}��F3t+D�e�]��\��ˋ|��yT�E�G�����[�t�<x�y)�<�C���z�O�ˡ]�ӯA�̓�-yʩ@M��LB�Y����Q�]ۑ#��-p:�5��=�`T'r(�7��P�	VJr ���X���4�5��\�B���Z�#�0��K�L&�\<�TxEQ z�+f��E����K��_�����8N?a�̓g\�hg���̼���EXG˳I�g�#G�Zᦓ/������F���kMJ��lF�n�Bi3�m��(
��֏+^�?�uԲ�q��8�� �CD���Cq�
Q�?��_(����YȈo��&�����J��W�2��F�y�{2�4x,���]�uh�]�������*��bY�3�RTtj���-�4�R��d�)�n��q�����[�;��hӠ�ڇ>í?	�]� ,��_p���hկy�v�p	m�l�D���,�"/���F���'΅Oo�'<��˰6ok��r���⒨���C!�pg�~WO���b(��<�y+VO<;1�Y��$~���C6@ef�s�:�?��m9�}��085�l}�=���GaS�^��ZX	>a�xx�ڿ��p@�x��?s�7�IL��~�%�w��E}|����_T�@8')��W���;��h��������H���(�oM-��*a�7$���j�ϝ>Pҧ�%<�Ccuۈ/W���ڷ��W��c+:L�=���ܯx����۟����MK���ԁ'��Ac��+a'�_NT�}Rx���YP,��r7ö��!���O���'.���Q�8�� #�O���X���wd^}�xW��K�ߝDm�N���Vb� W�اz7h)�TCEg(�hf\�QY�k��bR߂���_T���+Kx1�Dt�N5��R��́Ǵ(���u_���7��~N2�;�3P?�MpB� �=�ħr�po�!�D�c�R�]�3��mU�qڤ�A5A͜D"�T,{��D��ص�v�X���������?F0�]�r�ɓŇLBP� 
�Q��1/iC�OGGp��@Jl<�û���/��/w�`��5�����1��j�ZL�&{3,ݾ����͏qn����?�b�a�'/��=�	�����]�����p�aH�۩xW���?��i;Ol�JF�q��憇�Q�1���!��`������8A�*p;����B�1n&����cH�@z�kP�uGy&*�/n~�����h!�㹾�4~s��p���ܸ=uK�B�)���=��/��+�;?~l�f�i�jX���A1Hf��G����'J7� ��t�i�@�e�a���"�� �����S�R.�������9��Q`lL��]8�]����u�F��g����}l=�(��+��~{���1�#0[hO
���7����mPX~���a����mSmRJ��
��;�\U���S������}>�%m7����%>��>����IN��ɑR��g����U�Z\�XD����/�/����ޏ���H��ar�h���g�o���\�f�>	>�韐���N��@�_=��S�l�28�⌔5%�e'e��S��J�^��"(o�bb׿�4�[�\�>rEy��dhv6w��3���:o����j{Ĳ�z#���^��p,�ԩ�lB2LɄ[�� ?��]�^r7G,ͯ�����f&����p�+y�.�[䗐)�p�28�廡���-?n<�|��\���`;ꘕ�qB�Cn�E���ґ��]�Xӈ�W?�{�UGNM�6��p�ؙp"�QS�H�{	� �w�{��C�����w������z+�%y����[��(�6��6�m��@\�-3��]	/95�վiH2z>��Q!�d�62+��AK$..=��3��BQ�}�r/l"#��x�r�r����w��S��O4�z�eHL��"=��n܃&�.��3�6�h�k�aK�渓ٛ���P��a&�h�hg���hL;��;E��+����&;i^�#��kBD��J_�Z���;x=m��}��aS.�f�$z(t?��0���A�0���ݶ۬��&������y�f�ݯ¬gn�]��SE
�GL����f�.7Z��5")#��x))� �HDL
�������l��0x��?�D��X����8�H왣�����k���`h��B�Q�`��o��䓭?���M0������Ϲ�bw��89��L�K�ZA�����l|H��o!E'_�������\�W_���磈I��`ְy�E;Wv�jANJG%~'*g�����yP}ڼ<-k D��Ϫ�khS��
�VN�ہ��<j��v4 6 Qhn�4����}(�:ܵ��t:�C��oػ��b܈g�	n��w��xDB1�ȭ(�fA؊��PD��zG��׾\���[�mbgX���������QP�=��{A�uaH��#����2d<M?�l��e�����$���r�=7dHE"��9��'�K�>�K(r�g�P���rm>��2��f� ���B���d�;*B񔬪O���;��X�J遑���z3��Zc{$
"nK(o��K"���"���s"�����d|�ˏ������&+	I���"�Z���襡��qIP�w��%�0^���r��� E~���&K�����	¯Q����Fm�Ҁ�L8����pf�fR��S�-��F�{��B:�?8�o"_c�'g��_� {�c%�m%g�u�xM�A��$�����bU� �"	Ǡ(�܇�^�9�����%.�K@�k���<!.���_a.�:���hj��uɈp���Y�a�n��.pS�|�fW��%�JPD�L�5˾�uh(�Y�C½ ���zLZ���4[����ٞ$�y,+�$��i4yI�>��]�1�i��X��D��e8�U�ó�s����n�J�_��[t|5/ZWWͺ^��^4���24w)��vg���M�ͧo�ؾ�o@s�S�����9g�Dx��x���$�܀.W�*Ų�!�`:%�hډ?�������:��*���{o����WX$	VIT$VE��V0��kx�OYWAE�
��	3�r�!͐&�t�����힞��a�}�������U�:��9UNm�zmq��!Z��מ��W�X�V�y}w��-���J�%����҈n���?�ǧU5Ț�CۃZ��@����4�ۃwr��'�H��j5�.V�����J˙=��mRB
���X�p�i�p����HCs�x�-Ըn#y�?���r�e��"�y����#t�+�Q-�����7�X���k�|� �V�˪��s���^Щ�}��J<���\�/?�"���\��Ѵ�&I
~ⶡT��q59n|��/n�ﻼ��Ԑ���;
����^���gz�)(_�1�u���Nۥ?���/̥6��ҭo�55<�*�r��ך�s����8%�@�i���h��B�o��nq �sҖнzJ�ǱW�l�N�r� �-L��ǵs~����osdcQVֶ�s��zQC�5n�A6�:�e�Ay[��2_]L��;�3K�[��h%_�D�"��J��P�_��x�$�5[�5-Yf�K�!`!L�SW&=���^_>CM/~�� �_Á	�.N�<�z��u$;�3�)���,�a�l<�G����6�Fӂ��Z%#ːZ`llqHV��^�,l�r�Fy>�|���@V��n ���	�6q�<+1O#�F8�9l�&2B-~ ��c�ð�RU�-D�/+o�1��#]�̂دUahP7kV[��a7����-.�-`a�>��9A�@��j��()Р�ff���Ec��:_ۆo�6�x �j2D��*3�PEv���e��4�BG�[�@c��6�!䊥:F�������$C�L��U��t�DJ�X|U��;F��+�Y\���B�q#�Ζ�LJ�@ʒm��m�=�޺/�8#-R  <���c�*5vN�����X1�V䆊K�4$��̫ߣ�A��r�S���0�}��o�>>� 7 !�*�6�A;A��@L�+Qްc�\FSM�}G�h@�[H��ւ����$;个%�ޠ�s�J ��Z �0����KӇM�m��#R*��ߓw�� ������0/���[�<��T���HL�_hO(Y������*��NE��,��;�z݃���^��b�
�����P-�����`�{N�7W}
u����h�����s ���A��ؐ�<�#y��[�C���=���@�&&jE�0�P�_��(�3s
�^~�I�w��U�g��#�8=���缞eum�_��vVp0¡(�5���ڏ��Z��V���m��)�b[�O�0�xi���a��פ.;���e3�YjC)��=�MX�O�|t��[���������kgJ�����Dȣ<+5"6.���;��>p<��g��5BFWuO�#�� !��q�.v�6FFv}����0Ya����n�L���z��{0��;~ܡg|�m��^g�����$��-;J��U�y_LY���I()�1>�7�yz��8il�<G���`�rF.�zpcV�d�:�;8��٤��]�77m'���&�O�PF�'�f���L��8~x��bԂ�ߨ9%c�r}��]�n�*��CF���z��*�&�	�#�l�V���1ӵ"ݿ6VQ����)?��T���ke�f9�2��*�������~W�>������
ĳШ82��z�V��p�|�J=�5*a�(s��X����h͎t�E���<���r�s��+��Yf�v;UGu[,��B@ۨ���h,��*�=�vE�N�L�f�]ɺ涬��N��{��W����Vf�P�����c�x�ڕψ�]�Z�3xx�d����˺z5�1��J��F��D�u ��oL���� ���%\CR0��[���ƶƤ%�h��4SI��0Z�:Y�Fe[�?F�Ι�ZK�Le�Xx)pt�^�V�ӣ�=E��=�^��_f"�U�K��y�����LD�W� %�,h���?|����m��h���s��s������N�7�%���5_�|v7gu]��5��OӰ[��彄'�@B%�ʍ9-b�]�q(LC�ܯ��%�a!�*�/Cj��^o��^�0|��Y`W�資�&eրv��c��KcO{	�w�-m�~b�[P�KL�J��ʠ7�`�*�T����/�#U��������Nҭ�:˿�r��:����٠�;��8��6���ޘ��/n�*���}���I�J��5��^ӂ��&)^/=е�<}�Q���<g�s������W~J3ҿ��CE� F�	�|�!?�v���h��҂`�XT��	�ٍr���v����/�A�����+˔��هaD�C�fH��D�C{T��ٜ҆�S��Uf�|cU� Զ�]م�*"E�� [�����]c�]T��{+!��6 �c\2�#5^0+/���T� -^��f�3 � l�t��z6��9cǨ���aH�7�|2,3�~�e��O�qX��F�Jb68Q��|�5�̎lH�����^��?;�o���	����/t�"�(��.�#1��ͅ�ޯ�݅��k���p�����4`��KQ��-�n:�����Z��Q����V���@{)/����6���N����rK�/�(S�ŊQs!.�B�"���8�=��T�<�Zպr�S vL�X'�� $Ef7Ya�3���ѹP�A�.�h���z�ə4g�c���y���(3���q:����	:����K*�;��-L��2`�2�U�~6'�j�<k�+2؁ca�E@0,��:�Qv��J��뗝�Ȉ�	����&�~���S��\WA�b"&��f�Z6���?3g��o��f�5!����T�'��p���E�����v�]���f+�N�5{�����0�x�&v-��K�������F�o���[bH>VG��6n)�����;�X<t�2�������F!��d�;AC:���k���Ky��A�t�L��^Gϟ��|�M�m̭�4��j]�Gv��.�����v'MM����2"�`ưkhw���#B�kF/�qh7M����P>���(��1��eq�{�,�mzi��<jU�'w	��g�ejj��K3�z�+7=�0�rEX�c���p��u3d禯�k��f'Sؠ�s4
�ز[����[�V\���M�k����.r�_PY����?4���u��)X�{m-?�Ы�__J��'�ve�*"���%�4�t&u�O霢�:�T��9��?H[�u��7�2�2�$����7#s�1&����_q��x1~�Bԯ���yt��I�V�9 'K���cE�#V^z�pХ���=O��Ri�Ayv͗��g3�<�I�M�q��8����S���Q�6n�˭������s83`�z��C����d:��V$6̉	�swV�EV��"�F���^�~�Ըv2t�������.|bS�T�1|S^X��n�Х���хo+q��|���~xGl���۳Q�:�dp6˄�K�$r�� ��{6��-n���l<~>[:��Ә~����+�	=��\� �2�����4�ګ)F[�n
^��`ˍS���K��j���G�������C0i�Dƒy1C�P��#�t��+V�ڌ5x^�ݟo.���c(�DD�# �g��-�4�T��r��,�eF�/�n���g��A� 9��3���^U��:�p�MŦ�H����cl�)ݚ2^Y�w;V�s�{�8�a�����K[��MA_������40¾-<���;���'�sx{hԆ����]]h]N�8��/6���6o��S�F^Z��Y��0 �29��#Y%�*�MeH���#��N�y��JN�� �^���v���a3z��I�ɖ���ed�&��Hw|dd��|�m]�T��&ޥ��=������ϳ�7����Ұ�Oq"����>Z�7�K��RO�ߑ'���썪�ǐ�R}&�9x�)Z�	,���-cos���T7��������[	�H���*��M8�e�9E�5M#V��W��˒�s�?�����S�����N'=ک����8�,c%0�B��r�x�9��(��s�`��5�q��Iu�� p��>"��_�5/���;�&Q���%���a�U��,�O2�\�h}�v�kNu㥥��I�͈���b�3�V��P9QW'��P�
{�(쒔�>|�:����c��<��q�*Q6�3J�-nw(�[x��M�v�L��#K�6�w�w�������3PG�6��qIg��1_%���{�m�W��Y(py���,�}	H�ß9c4�$���X0�20�ݝ\��ŷy�9]�؜�̀�i�M�\�|_?�i�gY���%���qΩ��X���]���p�ЙB�<��P�ImL6EYv��3ߴ����"9�#�1�T���8%���2ݺ~>ˉ1S�f�I�3f{Q~�g�t�F��b�[P����C ���|�ka'p�R�y|���J�S
��,�t�X�nO�]	X�����J zG���Y�9�V�Y)��yt}$���B6`į*Dޛ5�c���,��V(�wx�Z ޾���r��ssc�vU*֦O`-O`]F��������3��xԆc��(��a8��e�	`�!�`�}���ƪ�w�� R:&x>�}�dp�oʊ$U�a�A_x�w���0���J3`_��$���%���댦���;	�� '�E�=蠽g��gp�'�feyK7�x��G!c�S(�d�n��z*,��4Q����EQq�˰H\�J��K>����,<��>ʷ�Ernk�ة/�&� W1w����<��usc�_��$�J�D�k����I��aR�a�׮&q�4+�\"���F�AB$��A<h. ����
�euvz}V�RT;a�L�r�,�8 /^^㢙C�I�R0%A�-��u��z��SCo� ��QI�B/�t��:��L�x�$U�ߦ
���E�7����f�M�>@�����g�d�+�ۅx�R��gV�Q�ۋ�\ԣ�G�:�.���;7��-��8}�Xt�)��$�ky������W�/���4�@��K����>��3{I���S�� Sc�SQ����F6���B�YmK����������C����!�O;�'�#t@}��0ni<m=f�f�@�B|�9���'�gz�*�-s&�q%��FQZ� /NM�?��,� ���b�[���[�@s��Ν	K���V��o�uIXTP��o �qu���N���.� �q�q����e��bwiEߊ��x��\l�u�tG*�l�}zy���_o/�ډ�媦2U� ���o���ݎ�-t3l<U����e�礱?U�ˠy�b��*�v�jq��%�HV�х<�^�1���[n��Ɖ��P߁��#�Vo��ޖ�
o����-��'ص��fsU��$�]��{�4�m)��WN~l�̋*�p�NK�8��H�
�5�ɀ�-{H�CE��֧��'>�`V�ٿ��a5��{�;�zP7���CMS8e���UZ�i�E���uA�|]����*~˸�"�A/����H��dЪr�U��K�^Ko�c���h|������G�3�����K����Рz���F�\��>���n"��`*��}N�|��*�
����|�%`���9D��Qe�F'����l�oV1�Ӣ�+R�G��e7�Q�]8}�9ߙ��0�x����nu�1�>�
��Jgs��g��<UV@՟Մz'�B�+2�+~��z�0�RQ��7١��U�&;{?QP��F0.�ժDM�[^��G9,�]�ll�k�(�ԥs!�+]XШ�����x���!���!     IEND�B`�PK   �M�Z�M/��  m     jsons/user_defined.jsonŘ�o�6 �����q��|˒���.�j�TU��
aUU��>����Q�E�ċ�cll~/�Ṑ�ҩ+Y�E2N29s�YVI��pH��)Z9˿_��+�\�ů�@����s���\�����gUܹL�2��P�i*K�v~�m:�2��JΝDm:1]	a ����b�)���e���Z��UX&šm��j��0�!E1@" ��^�](&(������u�c����Q�d�r�hY�wR$�6�sg��d�~�TE�?��T���.0n�=�S_����s���n���V�˶��P&����)�WIs�I��p��D08G���pU��Ze�C^���塬U��~ �T�3�|�� �m �7 tC򖀵l ���G��@������ZB#LK`��A� p-���8� �a `��v�wH�����xZ=-�3 #��1ϒ�J�rg��^�3��`��{Do���Fz���{D�5��{�Έ�#x�QtB/6:cv�`6c�7�Q�G��A��Fg���f,�n�3r�l3z����1����v#��C��r��bB/7�-&u6L�C�Ť��z��Po1��z���o1�>��^"Xo8.&��^q<T\Lz�c��x踘43a��x(��4���Ĥ��B��E'F�m�;Do:1�n�l#��Iu��'ѻNL�[-��^vb���[��m'&ۭ>i�^wb����L�;1�n��I�����g�H�O��4ab�z���w:	���mg��Y!�����k�=%���)ʼ��!鲠.@��̝���E��H~Z7{�5��d���F5�ӧl��W~�
�$U���X)�#�z4w��Y��.e���6�z��$̳6`�c�r����BL�J	<E��c&��)T�<���O֐�i��ˋ<�� +U��]��8�?�l��/�}�����z�k)�oy}�����k�aJݎ��:3�m<@�<^�p�� �؍��傍��<�dP$�PI0�@캄3�X�]o�L�/D�Bdj�u�P�Ej�k�T)x~�c��[_|P�X�j�?Y�۬>�6[�X[3n6�P�X�������d}���u�����"S;!�H���_Wk�L�D�7�YY�j����d�![�jգ�G�gl��e���ӈm�۫��:��vQ���cN�g����<�B�#O�g�B 1�,�=N=6y>���/PK
   �M�Z�
Bv;	  �I                   cirkitFile.jsonPK
   �M�Z��'S4  N4  /             h	  images/90a7334e-e219-40c9-b800-02625da96495.pngPK
   �M�Z��?�� � /             >  images/935ecb41-e360-41de-b535-f88365900f7a.pngPK
   �M�Zr�>�� � /             .D images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.pngPK
   �M�Z?��O�o  �o  /             :' images/ffe61187-e64a-4024-8cee-95dd034d2257.pngPK
   �M�Z�M/��  m               t� jsons/user_defined.jsonPK      �  j�   